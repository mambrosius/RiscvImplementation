`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module InstructionMemory(
  input         clock,
  input  [31:0] io_pc,
  output [31:0] io_inst
);
  reg [7:0] rom [0:239];
  reg [31:0] _GEN_0;
  wire [7:0] rom__T_790_data;
  wire [7:0] rom__T_790_addr;
  reg [31:0] _GEN_1;
  wire [7:0] rom__T_795_data;
  wire [7:0] rom__T_795_addr;
  reg [31:0] _GEN_2;
  wire [7:0] rom__T_800_data;
  wire [7:0] rom__T_800_addr;
  reg [31:0] _GEN_3;
  wire [7:0] rom__T_802_data;
  wire [7:0] rom__T_802_addr;
  reg [31:0] _GEN_4;
  wire [7:0] rom__T_8_data;
  wire [7:0] rom__T_8_addr;
  wire  rom__T_8_mask;
  wire  rom__T_8_en;
  wire [7:0] rom__T_11_data;
  wire [7:0] rom__T_11_addr;
  wire  rom__T_11_mask;
  wire  rom__T_11_en;
  wire [7:0] rom__T_14_data;
  wire [7:0] rom__T_14_addr;
  wire  rom__T_14_mask;
  wire  rom__T_14_en;
  wire [7:0] rom__T_17_data;
  wire [7:0] rom__T_17_addr;
  wire  rom__T_17_mask;
  wire  rom__T_17_en;
  wire [7:0] rom__T_21_data;
  wire [7:0] rom__T_21_addr;
  wire  rom__T_21_mask;
  wire  rom__T_21_en;
  wire [7:0] rom__T_24_data;
  wire [7:0] rom__T_24_addr;
  wire  rom__T_24_mask;
  wire  rom__T_24_en;
  wire [7:0] rom__T_27_data;
  wire [7:0] rom__T_27_addr;
  wire  rom__T_27_mask;
  wire  rom__T_27_en;
  wire [7:0] rom__T_30_data;
  wire [7:0] rom__T_30_addr;
  wire  rom__T_30_mask;
  wire  rom__T_30_en;
  wire [7:0] rom__T_34_data;
  wire [7:0] rom__T_34_addr;
  wire  rom__T_34_mask;
  wire  rom__T_34_en;
  wire [7:0] rom__T_37_data;
  wire [7:0] rom__T_37_addr;
  wire  rom__T_37_mask;
  wire  rom__T_37_en;
  wire [7:0] rom__T_40_data;
  wire [7:0] rom__T_40_addr;
  wire  rom__T_40_mask;
  wire  rom__T_40_en;
  wire [7:0] rom__T_43_data;
  wire [7:0] rom__T_43_addr;
  wire  rom__T_43_mask;
  wire  rom__T_43_en;
  wire [7:0] rom__T_47_data;
  wire [7:0] rom__T_47_addr;
  wire  rom__T_47_mask;
  wire  rom__T_47_en;
  wire [7:0] rom__T_50_data;
  wire [7:0] rom__T_50_addr;
  wire  rom__T_50_mask;
  wire  rom__T_50_en;
  wire [7:0] rom__T_53_data;
  wire [7:0] rom__T_53_addr;
  wire  rom__T_53_mask;
  wire  rom__T_53_en;
  wire [7:0] rom__T_56_data;
  wire [7:0] rom__T_56_addr;
  wire  rom__T_56_mask;
  wire  rom__T_56_en;
  wire [7:0] rom__T_60_data;
  wire [7:0] rom__T_60_addr;
  wire  rom__T_60_mask;
  wire  rom__T_60_en;
  wire [7:0] rom__T_63_data;
  wire [7:0] rom__T_63_addr;
  wire  rom__T_63_mask;
  wire  rom__T_63_en;
  wire [7:0] rom__T_66_data;
  wire [7:0] rom__T_66_addr;
  wire  rom__T_66_mask;
  wire  rom__T_66_en;
  wire [7:0] rom__T_69_data;
  wire [7:0] rom__T_69_addr;
  wire  rom__T_69_mask;
  wire  rom__T_69_en;
  wire [7:0] rom__T_73_data;
  wire [7:0] rom__T_73_addr;
  wire  rom__T_73_mask;
  wire  rom__T_73_en;
  wire [7:0] rom__T_76_data;
  wire [7:0] rom__T_76_addr;
  wire  rom__T_76_mask;
  wire  rom__T_76_en;
  wire [7:0] rom__T_79_data;
  wire [7:0] rom__T_79_addr;
  wire  rom__T_79_mask;
  wire  rom__T_79_en;
  wire [7:0] rom__T_82_data;
  wire [7:0] rom__T_82_addr;
  wire  rom__T_82_mask;
  wire  rom__T_82_en;
  wire [7:0] rom__T_86_data;
  wire [7:0] rom__T_86_addr;
  wire  rom__T_86_mask;
  wire  rom__T_86_en;
  wire [7:0] rom__T_89_data;
  wire [7:0] rom__T_89_addr;
  wire  rom__T_89_mask;
  wire  rom__T_89_en;
  wire [7:0] rom__T_92_data;
  wire [7:0] rom__T_92_addr;
  wire  rom__T_92_mask;
  wire  rom__T_92_en;
  wire [7:0] rom__T_95_data;
  wire [7:0] rom__T_95_addr;
  wire  rom__T_95_mask;
  wire  rom__T_95_en;
  wire [7:0] rom__T_99_data;
  wire [7:0] rom__T_99_addr;
  wire  rom__T_99_mask;
  wire  rom__T_99_en;
  wire [7:0] rom__T_102_data;
  wire [7:0] rom__T_102_addr;
  wire  rom__T_102_mask;
  wire  rom__T_102_en;
  wire [7:0] rom__T_105_data;
  wire [7:0] rom__T_105_addr;
  wire  rom__T_105_mask;
  wire  rom__T_105_en;
  wire [7:0] rom__T_108_data;
  wire [7:0] rom__T_108_addr;
  wire  rom__T_108_mask;
  wire  rom__T_108_en;
  wire [7:0] rom__T_112_data;
  wire [7:0] rom__T_112_addr;
  wire  rom__T_112_mask;
  wire  rom__T_112_en;
  wire [7:0] rom__T_115_data;
  wire [7:0] rom__T_115_addr;
  wire  rom__T_115_mask;
  wire  rom__T_115_en;
  wire [7:0] rom__T_118_data;
  wire [7:0] rom__T_118_addr;
  wire  rom__T_118_mask;
  wire  rom__T_118_en;
  wire [7:0] rom__T_121_data;
  wire [7:0] rom__T_121_addr;
  wire  rom__T_121_mask;
  wire  rom__T_121_en;
  wire [7:0] rom__T_125_data;
  wire [7:0] rom__T_125_addr;
  wire  rom__T_125_mask;
  wire  rom__T_125_en;
  wire [7:0] rom__T_128_data;
  wire [7:0] rom__T_128_addr;
  wire  rom__T_128_mask;
  wire  rom__T_128_en;
  wire [7:0] rom__T_131_data;
  wire [7:0] rom__T_131_addr;
  wire  rom__T_131_mask;
  wire  rom__T_131_en;
  wire [7:0] rom__T_134_data;
  wire [7:0] rom__T_134_addr;
  wire  rom__T_134_mask;
  wire  rom__T_134_en;
  wire [7:0] rom__T_138_data;
  wire [7:0] rom__T_138_addr;
  wire  rom__T_138_mask;
  wire  rom__T_138_en;
  wire [7:0] rom__T_141_data;
  wire [7:0] rom__T_141_addr;
  wire  rom__T_141_mask;
  wire  rom__T_141_en;
  wire [7:0] rom__T_144_data;
  wire [7:0] rom__T_144_addr;
  wire  rom__T_144_mask;
  wire  rom__T_144_en;
  wire [7:0] rom__T_147_data;
  wire [7:0] rom__T_147_addr;
  wire  rom__T_147_mask;
  wire  rom__T_147_en;
  wire [7:0] rom__T_151_data;
  wire [7:0] rom__T_151_addr;
  wire  rom__T_151_mask;
  wire  rom__T_151_en;
  wire [7:0] rom__T_154_data;
  wire [7:0] rom__T_154_addr;
  wire  rom__T_154_mask;
  wire  rom__T_154_en;
  wire [7:0] rom__T_157_data;
  wire [7:0] rom__T_157_addr;
  wire  rom__T_157_mask;
  wire  rom__T_157_en;
  wire [7:0] rom__T_160_data;
  wire [7:0] rom__T_160_addr;
  wire  rom__T_160_mask;
  wire  rom__T_160_en;
  wire [7:0] rom__T_164_data;
  wire [7:0] rom__T_164_addr;
  wire  rom__T_164_mask;
  wire  rom__T_164_en;
  wire [7:0] rom__T_167_data;
  wire [7:0] rom__T_167_addr;
  wire  rom__T_167_mask;
  wire  rom__T_167_en;
  wire [7:0] rom__T_170_data;
  wire [7:0] rom__T_170_addr;
  wire  rom__T_170_mask;
  wire  rom__T_170_en;
  wire [7:0] rom__T_173_data;
  wire [7:0] rom__T_173_addr;
  wire  rom__T_173_mask;
  wire  rom__T_173_en;
  wire [7:0] rom__T_177_data;
  wire [7:0] rom__T_177_addr;
  wire  rom__T_177_mask;
  wire  rom__T_177_en;
  wire [7:0] rom__T_180_data;
  wire [7:0] rom__T_180_addr;
  wire  rom__T_180_mask;
  wire  rom__T_180_en;
  wire [7:0] rom__T_183_data;
  wire [7:0] rom__T_183_addr;
  wire  rom__T_183_mask;
  wire  rom__T_183_en;
  wire [7:0] rom__T_186_data;
  wire [7:0] rom__T_186_addr;
  wire  rom__T_186_mask;
  wire  rom__T_186_en;
  wire [7:0] rom__T_190_data;
  wire [7:0] rom__T_190_addr;
  wire  rom__T_190_mask;
  wire  rom__T_190_en;
  wire [7:0] rom__T_193_data;
  wire [7:0] rom__T_193_addr;
  wire  rom__T_193_mask;
  wire  rom__T_193_en;
  wire [7:0] rom__T_196_data;
  wire [7:0] rom__T_196_addr;
  wire  rom__T_196_mask;
  wire  rom__T_196_en;
  wire [7:0] rom__T_199_data;
  wire [7:0] rom__T_199_addr;
  wire  rom__T_199_mask;
  wire  rom__T_199_en;
  wire [7:0] rom__T_203_data;
  wire [7:0] rom__T_203_addr;
  wire  rom__T_203_mask;
  wire  rom__T_203_en;
  wire [7:0] rom__T_206_data;
  wire [7:0] rom__T_206_addr;
  wire  rom__T_206_mask;
  wire  rom__T_206_en;
  wire [7:0] rom__T_209_data;
  wire [7:0] rom__T_209_addr;
  wire  rom__T_209_mask;
  wire  rom__T_209_en;
  wire [7:0] rom__T_212_data;
  wire [7:0] rom__T_212_addr;
  wire  rom__T_212_mask;
  wire  rom__T_212_en;
  wire [7:0] rom__T_216_data;
  wire [7:0] rom__T_216_addr;
  wire  rom__T_216_mask;
  wire  rom__T_216_en;
  wire [7:0] rom__T_219_data;
  wire [7:0] rom__T_219_addr;
  wire  rom__T_219_mask;
  wire  rom__T_219_en;
  wire [7:0] rom__T_222_data;
  wire [7:0] rom__T_222_addr;
  wire  rom__T_222_mask;
  wire  rom__T_222_en;
  wire [7:0] rom__T_225_data;
  wire [7:0] rom__T_225_addr;
  wire  rom__T_225_mask;
  wire  rom__T_225_en;
  wire [7:0] rom__T_229_data;
  wire [7:0] rom__T_229_addr;
  wire  rom__T_229_mask;
  wire  rom__T_229_en;
  wire [7:0] rom__T_232_data;
  wire [7:0] rom__T_232_addr;
  wire  rom__T_232_mask;
  wire  rom__T_232_en;
  wire [7:0] rom__T_235_data;
  wire [7:0] rom__T_235_addr;
  wire  rom__T_235_mask;
  wire  rom__T_235_en;
  wire [7:0] rom__T_238_data;
  wire [7:0] rom__T_238_addr;
  wire  rom__T_238_mask;
  wire  rom__T_238_en;
  wire [7:0] rom__T_242_data;
  wire [7:0] rom__T_242_addr;
  wire  rom__T_242_mask;
  wire  rom__T_242_en;
  wire [7:0] rom__T_245_data;
  wire [7:0] rom__T_245_addr;
  wire  rom__T_245_mask;
  wire  rom__T_245_en;
  wire [7:0] rom__T_248_data;
  wire [7:0] rom__T_248_addr;
  wire  rom__T_248_mask;
  wire  rom__T_248_en;
  wire [7:0] rom__T_251_data;
  wire [7:0] rom__T_251_addr;
  wire  rom__T_251_mask;
  wire  rom__T_251_en;
  wire [7:0] rom__T_255_data;
  wire [7:0] rom__T_255_addr;
  wire  rom__T_255_mask;
  wire  rom__T_255_en;
  wire [7:0] rom__T_258_data;
  wire [7:0] rom__T_258_addr;
  wire  rom__T_258_mask;
  wire  rom__T_258_en;
  wire [7:0] rom__T_261_data;
  wire [7:0] rom__T_261_addr;
  wire  rom__T_261_mask;
  wire  rom__T_261_en;
  wire [7:0] rom__T_264_data;
  wire [7:0] rom__T_264_addr;
  wire  rom__T_264_mask;
  wire  rom__T_264_en;
  wire [7:0] rom__T_268_data;
  wire [7:0] rom__T_268_addr;
  wire  rom__T_268_mask;
  wire  rom__T_268_en;
  wire [7:0] rom__T_271_data;
  wire [7:0] rom__T_271_addr;
  wire  rom__T_271_mask;
  wire  rom__T_271_en;
  wire [7:0] rom__T_274_data;
  wire [7:0] rom__T_274_addr;
  wire  rom__T_274_mask;
  wire  rom__T_274_en;
  wire [7:0] rom__T_277_data;
  wire [7:0] rom__T_277_addr;
  wire  rom__T_277_mask;
  wire  rom__T_277_en;
  wire [7:0] rom__T_281_data;
  wire [7:0] rom__T_281_addr;
  wire  rom__T_281_mask;
  wire  rom__T_281_en;
  wire [7:0] rom__T_284_data;
  wire [7:0] rom__T_284_addr;
  wire  rom__T_284_mask;
  wire  rom__T_284_en;
  wire [7:0] rom__T_287_data;
  wire [7:0] rom__T_287_addr;
  wire  rom__T_287_mask;
  wire  rom__T_287_en;
  wire [7:0] rom__T_290_data;
  wire [7:0] rom__T_290_addr;
  wire  rom__T_290_mask;
  wire  rom__T_290_en;
  wire [7:0] rom__T_294_data;
  wire [7:0] rom__T_294_addr;
  wire  rom__T_294_mask;
  wire  rom__T_294_en;
  wire [7:0] rom__T_297_data;
  wire [7:0] rom__T_297_addr;
  wire  rom__T_297_mask;
  wire  rom__T_297_en;
  wire [7:0] rom__T_300_data;
  wire [7:0] rom__T_300_addr;
  wire  rom__T_300_mask;
  wire  rom__T_300_en;
  wire [7:0] rom__T_303_data;
  wire [7:0] rom__T_303_addr;
  wire  rom__T_303_mask;
  wire  rom__T_303_en;
  wire [7:0] rom__T_307_data;
  wire [7:0] rom__T_307_addr;
  wire  rom__T_307_mask;
  wire  rom__T_307_en;
  wire [7:0] rom__T_310_data;
  wire [7:0] rom__T_310_addr;
  wire  rom__T_310_mask;
  wire  rom__T_310_en;
  wire [7:0] rom__T_313_data;
  wire [7:0] rom__T_313_addr;
  wire  rom__T_313_mask;
  wire  rom__T_313_en;
  wire [7:0] rom__T_316_data;
  wire [7:0] rom__T_316_addr;
  wire  rom__T_316_mask;
  wire  rom__T_316_en;
  wire [7:0] rom__T_320_data;
  wire [7:0] rom__T_320_addr;
  wire  rom__T_320_mask;
  wire  rom__T_320_en;
  wire [7:0] rom__T_323_data;
  wire [7:0] rom__T_323_addr;
  wire  rom__T_323_mask;
  wire  rom__T_323_en;
  wire [7:0] rom__T_326_data;
  wire [7:0] rom__T_326_addr;
  wire  rom__T_326_mask;
  wire  rom__T_326_en;
  wire [7:0] rom__T_329_data;
  wire [7:0] rom__T_329_addr;
  wire  rom__T_329_mask;
  wire  rom__T_329_en;
  wire [7:0] rom__T_333_data;
  wire [7:0] rom__T_333_addr;
  wire  rom__T_333_mask;
  wire  rom__T_333_en;
  wire [7:0] rom__T_336_data;
  wire [7:0] rom__T_336_addr;
  wire  rom__T_336_mask;
  wire  rom__T_336_en;
  wire [7:0] rom__T_339_data;
  wire [7:0] rom__T_339_addr;
  wire  rom__T_339_mask;
  wire  rom__T_339_en;
  wire [7:0] rom__T_342_data;
  wire [7:0] rom__T_342_addr;
  wire  rom__T_342_mask;
  wire  rom__T_342_en;
  wire [7:0] rom__T_346_data;
  wire [7:0] rom__T_346_addr;
  wire  rom__T_346_mask;
  wire  rom__T_346_en;
  wire [7:0] rom__T_349_data;
  wire [7:0] rom__T_349_addr;
  wire  rom__T_349_mask;
  wire  rom__T_349_en;
  wire [7:0] rom__T_352_data;
  wire [7:0] rom__T_352_addr;
  wire  rom__T_352_mask;
  wire  rom__T_352_en;
  wire [7:0] rom__T_355_data;
  wire [7:0] rom__T_355_addr;
  wire  rom__T_355_mask;
  wire  rom__T_355_en;
  wire [7:0] rom__T_359_data;
  wire [7:0] rom__T_359_addr;
  wire  rom__T_359_mask;
  wire  rom__T_359_en;
  wire [7:0] rom__T_362_data;
  wire [7:0] rom__T_362_addr;
  wire  rom__T_362_mask;
  wire  rom__T_362_en;
  wire [7:0] rom__T_365_data;
  wire [7:0] rom__T_365_addr;
  wire  rom__T_365_mask;
  wire  rom__T_365_en;
  wire [7:0] rom__T_368_data;
  wire [7:0] rom__T_368_addr;
  wire  rom__T_368_mask;
  wire  rom__T_368_en;
  wire [7:0] rom__T_372_data;
  wire [7:0] rom__T_372_addr;
  wire  rom__T_372_mask;
  wire  rom__T_372_en;
  wire [7:0] rom__T_375_data;
  wire [7:0] rom__T_375_addr;
  wire  rom__T_375_mask;
  wire  rom__T_375_en;
  wire [7:0] rom__T_378_data;
  wire [7:0] rom__T_378_addr;
  wire  rom__T_378_mask;
  wire  rom__T_378_en;
  wire [7:0] rom__T_381_data;
  wire [7:0] rom__T_381_addr;
  wire  rom__T_381_mask;
  wire  rom__T_381_en;
  wire [7:0] rom__T_385_data;
  wire [7:0] rom__T_385_addr;
  wire  rom__T_385_mask;
  wire  rom__T_385_en;
  wire [7:0] rom__T_388_data;
  wire [7:0] rom__T_388_addr;
  wire  rom__T_388_mask;
  wire  rom__T_388_en;
  wire [7:0] rom__T_391_data;
  wire [7:0] rom__T_391_addr;
  wire  rom__T_391_mask;
  wire  rom__T_391_en;
  wire [7:0] rom__T_394_data;
  wire [7:0] rom__T_394_addr;
  wire  rom__T_394_mask;
  wire  rom__T_394_en;
  wire [7:0] rom__T_398_data;
  wire [7:0] rom__T_398_addr;
  wire  rom__T_398_mask;
  wire  rom__T_398_en;
  wire [7:0] rom__T_401_data;
  wire [7:0] rom__T_401_addr;
  wire  rom__T_401_mask;
  wire  rom__T_401_en;
  wire [7:0] rom__T_404_data;
  wire [7:0] rom__T_404_addr;
  wire  rom__T_404_mask;
  wire  rom__T_404_en;
  wire [7:0] rom__T_407_data;
  wire [7:0] rom__T_407_addr;
  wire  rom__T_407_mask;
  wire  rom__T_407_en;
  wire [7:0] rom__T_411_data;
  wire [7:0] rom__T_411_addr;
  wire  rom__T_411_mask;
  wire  rom__T_411_en;
  wire [7:0] rom__T_414_data;
  wire [7:0] rom__T_414_addr;
  wire  rom__T_414_mask;
  wire  rom__T_414_en;
  wire [7:0] rom__T_417_data;
  wire [7:0] rom__T_417_addr;
  wire  rom__T_417_mask;
  wire  rom__T_417_en;
  wire [7:0] rom__T_420_data;
  wire [7:0] rom__T_420_addr;
  wire  rom__T_420_mask;
  wire  rom__T_420_en;
  wire [7:0] rom__T_424_data;
  wire [7:0] rom__T_424_addr;
  wire  rom__T_424_mask;
  wire  rom__T_424_en;
  wire [7:0] rom__T_427_data;
  wire [7:0] rom__T_427_addr;
  wire  rom__T_427_mask;
  wire  rom__T_427_en;
  wire [7:0] rom__T_430_data;
  wire [7:0] rom__T_430_addr;
  wire  rom__T_430_mask;
  wire  rom__T_430_en;
  wire [7:0] rom__T_433_data;
  wire [7:0] rom__T_433_addr;
  wire  rom__T_433_mask;
  wire  rom__T_433_en;
  wire [7:0] rom__T_437_data;
  wire [7:0] rom__T_437_addr;
  wire  rom__T_437_mask;
  wire  rom__T_437_en;
  wire [7:0] rom__T_440_data;
  wire [7:0] rom__T_440_addr;
  wire  rom__T_440_mask;
  wire  rom__T_440_en;
  wire [7:0] rom__T_443_data;
  wire [7:0] rom__T_443_addr;
  wire  rom__T_443_mask;
  wire  rom__T_443_en;
  wire [7:0] rom__T_446_data;
  wire [7:0] rom__T_446_addr;
  wire  rom__T_446_mask;
  wire  rom__T_446_en;
  wire [7:0] rom__T_450_data;
  wire [7:0] rom__T_450_addr;
  wire  rom__T_450_mask;
  wire  rom__T_450_en;
  wire [7:0] rom__T_453_data;
  wire [7:0] rom__T_453_addr;
  wire  rom__T_453_mask;
  wire  rom__T_453_en;
  wire [7:0] rom__T_456_data;
  wire [7:0] rom__T_456_addr;
  wire  rom__T_456_mask;
  wire  rom__T_456_en;
  wire [7:0] rom__T_459_data;
  wire [7:0] rom__T_459_addr;
  wire  rom__T_459_mask;
  wire  rom__T_459_en;
  wire [7:0] rom__T_463_data;
  wire [7:0] rom__T_463_addr;
  wire  rom__T_463_mask;
  wire  rom__T_463_en;
  wire [7:0] rom__T_466_data;
  wire [7:0] rom__T_466_addr;
  wire  rom__T_466_mask;
  wire  rom__T_466_en;
  wire [7:0] rom__T_469_data;
  wire [7:0] rom__T_469_addr;
  wire  rom__T_469_mask;
  wire  rom__T_469_en;
  wire [7:0] rom__T_472_data;
  wire [7:0] rom__T_472_addr;
  wire  rom__T_472_mask;
  wire  rom__T_472_en;
  wire [7:0] rom__T_476_data;
  wire [7:0] rom__T_476_addr;
  wire  rom__T_476_mask;
  wire  rom__T_476_en;
  wire [7:0] rom__T_479_data;
  wire [7:0] rom__T_479_addr;
  wire  rom__T_479_mask;
  wire  rom__T_479_en;
  wire [7:0] rom__T_482_data;
  wire [7:0] rom__T_482_addr;
  wire  rom__T_482_mask;
  wire  rom__T_482_en;
  wire [7:0] rom__T_485_data;
  wire [7:0] rom__T_485_addr;
  wire  rom__T_485_mask;
  wire  rom__T_485_en;
  wire [7:0] rom__T_489_data;
  wire [7:0] rom__T_489_addr;
  wire  rom__T_489_mask;
  wire  rom__T_489_en;
  wire [7:0] rom__T_492_data;
  wire [7:0] rom__T_492_addr;
  wire  rom__T_492_mask;
  wire  rom__T_492_en;
  wire [7:0] rom__T_495_data;
  wire [7:0] rom__T_495_addr;
  wire  rom__T_495_mask;
  wire  rom__T_495_en;
  wire [7:0] rom__T_498_data;
  wire [7:0] rom__T_498_addr;
  wire  rom__T_498_mask;
  wire  rom__T_498_en;
  wire [7:0] rom__T_502_data;
  wire [7:0] rom__T_502_addr;
  wire  rom__T_502_mask;
  wire  rom__T_502_en;
  wire [7:0] rom__T_505_data;
  wire [7:0] rom__T_505_addr;
  wire  rom__T_505_mask;
  wire  rom__T_505_en;
  wire [7:0] rom__T_508_data;
  wire [7:0] rom__T_508_addr;
  wire  rom__T_508_mask;
  wire  rom__T_508_en;
  wire [7:0] rom__T_511_data;
  wire [7:0] rom__T_511_addr;
  wire  rom__T_511_mask;
  wire  rom__T_511_en;
  wire [7:0] rom__T_515_data;
  wire [7:0] rom__T_515_addr;
  wire  rom__T_515_mask;
  wire  rom__T_515_en;
  wire [7:0] rom__T_518_data;
  wire [7:0] rom__T_518_addr;
  wire  rom__T_518_mask;
  wire  rom__T_518_en;
  wire [7:0] rom__T_521_data;
  wire [7:0] rom__T_521_addr;
  wire  rom__T_521_mask;
  wire  rom__T_521_en;
  wire [7:0] rom__T_524_data;
  wire [7:0] rom__T_524_addr;
  wire  rom__T_524_mask;
  wire  rom__T_524_en;
  wire [7:0] rom__T_528_data;
  wire [7:0] rom__T_528_addr;
  wire  rom__T_528_mask;
  wire  rom__T_528_en;
  wire [7:0] rom__T_531_data;
  wire [7:0] rom__T_531_addr;
  wire  rom__T_531_mask;
  wire  rom__T_531_en;
  wire [7:0] rom__T_534_data;
  wire [7:0] rom__T_534_addr;
  wire  rom__T_534_mask;
  wire  rom__T_534_en;
  wire [7:0] rom__T_537_data;
  wire [7:0] rom__T_537_addr;
  wire  rom__T_537_mask;
  wire  rom__T_537_en;
  wire [7:0] rom__T_541_data;
  wire [7:0] rom__T_541_addr;
  wire  rom__T_541_mask;
  wire  rom__T_541_en;
  wire [7:0] rom__T_544_data;
  wire [7:0] rom__T_544_addr;
  wire  rom__T_544_mask;
  wire  rom__T_544_en;
  wire [7:0] rom__T_547_data;
  wire [7:0] rom__T_547_addr;
  wire  rom__T_547_mask;
  wire  rom__T_547_en;
  wire [7:0] rom__T_550_data;
  wire [7:0] rom__T_550_addr;
  wire  rom__T_550_mask;
  wire  rom__T_550_en;
  wire [7:0] rom__T_554_data;
  wire [7:0] rom__T_554_addr;
  wire  rom__T_554_mask;
  wire  rom__T_554_en;
  wire [7:0] rom__T_557_data;
  wire [7:0] rom__T_557_addr;
  wire  rom__T_557_mask;
  wire  rom__T_557_en;
  wire [7:0] rom__T_560_data;
  wire [7:0] rom__T_560_addr;
  wire  rom__T_560_mask;
  wire  rom__T_560_en;
  wire [7:0] rom__T_563_data;
  wire [7:0] rom__T_563_addr;
  wire  rom__T_563_mask;
  wire  rom__T_563_en;
  wire [7:0] rom__T_567_data;
  wire [7:0] rom__T_567_addr;
  wire  rom__T_567_mask;
  wire  rom__T_567_en;
  wire [7:0] rom__T_570_data;
  wire [7:0] rom__T_570_addr;
  wire  rom__T_570_mask;
  wire  rom__T_570_en;
  wire [7:0] rom__T_573_data;
  wire [7:0] rom__T_573_addr;
  wire  rom__T_573_mask;
  wire  rom__T_573_en;
  wire [7:0] rom__T_576_data;
  wire [7:0] rom__T_576_addr;
  wire  rom__T_576_mask;
  wire  rom__T_576_en;
  wire [7:0] rom__T_580_data;
  wire [7:0] rom__T_580_addr;
  wire  rom__T_580_mask;
  wire  rom__T_580_en;
  wire [7:0] rom__T_583_data;
  wire [7:0] rom__T_583_addr;
  wire  rom__T_583_mask;
  wire  rom__T_583_en;
  wire [7:0] rom__T_586_data;
  wire [7:0] rom__T_586_addr;
  wire  rom__T_586_mask;
  wire  rom__T_586_en;
  wire [7:0] rom__T_589_data;
  wire [7:0] rom__T_589_addr;
  wire  rom__T_589_mask;
  wire  rom__T_589_en;
  wire [7:0] rom__T_593_data;
  wire [7:0] rom__T_593_addr;
  wire  rom__T_593_mask;
  wire  rom__T_593_en;
  wire [7:0] rom__T_596_data;
  wire [7:0] rom__T_596_addr;
  wire  rom__T_596_mask;
  wire  rom__T_596_en;
  wire [7:0] rom__T_599_data;
  wire [7:0] rom__T_599_addr;
  wire  rom__T_599_mask;
  wire  rom__T_599_en;
  wire [7:0] rom__T_602_data;
  wire [7:0] rom__T_602_addr;
  wire  rom__T_602_mask;
  wire  rom__T_602_en;
  wire [7:0] rom__T_606_data;
  wire [7:0] rom__T_606_addr;
  wire  rom__T_606_mask;
  wire  rom__T_606_en;
  wire [7:0] rom__T_609_data;
  wire [7:0] rom__T_609_addr;
  wire  rom__T_609_mask;
  wire  rom__T_609_en;
  wire [7:0] rom__T_612_data;
  wire [7:0] rom__T_612_addr;
  wire  rom__T_612_mask;
  wire  rom__T_612_en;
  wire [7:0] rom__T_615_data;
  wire [7:0] rom__T_615_addr;
  wire  rom__T_615_mask;
  wire  rom__T_615_en;
  wire [7:0] rom__T_619_data;
  wire [7:0] rom__T_619_addr;
  wire  rom__T_619_mask;
  wire  rom__T_619_en;
  wire [7:0] rom__T_622_data;
  wire [7:0] rom__T_622_addr;
  wire  rom__T_622_mask;
  wire  rom__T_622_en;
  wire [7:0] rom__T_625_data;
  wire [7:0] rom__T_625_addr;
  wire  rom__T_625_mask;
  wire  rom__T_625_en;
  wire [7:0] rom__T_628_data;
  wire [7:0] rom__T_628_addr;
  wire  rom__T_628_mask;
  wire  rom__T_628_en;
  wire [7:0] rom__T_632_data;
  wire [7:0] rom__T_632_addr;
  wire  rom__T_632_mask;
  wire  rom__T_632_en;
  wire [7:0] rom__T_635_data;
  wire [7:0] rom__T_635_addr;
  wire  rom__T_635_mask;
  wire  rom__T_635_en;
  wire [7:0] rom__T_638_data;
  wire [7:0] rom__T_638_addr;
  wire  rom__T_638_mask;
  wire  rom__T_638_en;
  wire [7:0] rom__T_641_data;
  wire [7:0] rom__T_641_addr;
  wire  rom__T_641_mask;
  wire  rom__T_641_en;
  wire [7:0] rom__T_645_data;
  wire [7:0] rom__T_645_addr;
  wire  rom__T_645_mask;
  wire  rom__T_645_en;
  wire [7:0] rom__T_648_data;
  wire [7:0] rom__T_648_addr;
  wire  rom__T_648_mask;
  wire  rom__T_648_en;
  wire [7:0] rom__T_651_data;
  wire [7:0] rom__T_651_addr;
  wire  rom__T_651_mask;
  wire  rom__T_651_en;
  wire [7:0] rom__T_654_data;
  wire [7:0] rom__T_654_addr;
  wire  rom__T_654_mask;
  wire  rom__T_654_en;
  wire [7:0] rom__T_658_data;
  wire [7:0] rom__T_658_addr;
  wire  rom__T_658_mask;
  wire  rom__T_658_en;
  wire [7:0] rom__T_661_data;
  wire [7:0] rom__T_661_addr;
  wire  rom__T_661_mask;
  wire  rom__T_661_en;
  wire [7:0] rom__T_664_data;
  wire [7:0] rom__T_664_addr;
  wire  rom__T_664_mask;
  wire  rom__T_664_en;
  wire [7:0] rom__T_667_data;
  wire [7:0] rom__T_667_addr;
  wire  rom__T_667_mask;
  wire  rom__T_667_en;
  wire [7:0] rom__T_671_data;
  wire [7:0] rom__T_671_addr;
  wire  rom__T_671_mask;
  wire  rom__T_671_en;
  wire [7:0] rom__T_674_data;
  wire [7:0] rom__T_674_addr;
  wire  rom__T_674_mask;
  wire  rom__T_674_en;
  wire [7:0] rom__T_677_data;
  wire [7:0] rom__T_677_addr;
  wire  rom__T_677_mask;
  wire  rom__T_677_en;
  wire [7:0] rom__T_680_data;
  wire [7:0] rom__T_680_addr;
  wire  rom__T_680_mask;
  wire  rom__T_680_en;
  wire [7:0] rom__T_684_data;
  wire [7:0] rom__T_684_addr;
  wire  rom__T_684_mask;
  wire  rom__T_684_en;
  wire [7:0] rom__T_687_data;
  wire [7:0] rom__T_687_addr;
  wire  rom__T_687_mask;
  wire  rom__T_687_en;
  wire [7:0] rom__T_690_data;
  wire [7:0] rom__T_690_addr;
  wire  rom__T_690_mask;
  wire  rom__T_690_en;
  wire [7:0] rom__T_693_data;
  wire [7:0] rom__T_693_addr;
  wire  rom__T_693_mask;
  wire  rom__T_693_en;
  wire [7:0] rom__T_697_data;
  wire [7:0] rom__T_697_addr;
  wire  rom__T_697_mask;
  wire  rom__T_697_en;
  wire [7:0] rom__T_700_data;
  wire [7:0] rom__T_700_addr;
  wire  rom__T_700_mask;
  wire  rom__T_700_en;
  wire [7:0] rom__T_703_data;
  wire [7:0] rom__T_703_addr;
  wire  rom__T_703_mask;
  wire  rom__T_703_en;
  wire [7:0] rom__T_706_data;
  wire [7:0] rom__T_706_addr;
  wire  rom__T_706_mask;
  wire  rom__T_706_en;
  wire [7:0] rom__T_710_data;
  wire [7:0] rom__T_710_addr;
  wire  rom__T_710_mask;
  wire  rom__T_710_en;
  wire [7:0] rom__T_713_data;
  wire [7:0] rom__T_713_addr;
  wire  rom__T_713_mask;
  wire  rom__T_713_en;
  wire [7:0] rom__T_716_data;
  wire [7:0] rom__T_716_addr;
  wire  rom__T_716_mask;
  wire  rom__T_716_en;
  wire [7:0] rom__T_719_data;
  wire [7:0] rom__T_719_addr;
  wire  rom__T_719_mask;
  wire  rom__T_719_en;
  wire [7:0] rom__T_723_data;
  wire [7:0] rom__T_723_addr;
  wire  rom__T_723_mask;
  wire  rom__T_723_en;
  wire [7:0] rom__T_726_data;
  wire [7:0] rom__T_726_addr;
  wire  rom__T_726_mask;
  wire  rom__T_726_en;
  wire [7:0] rom__T_729_data;
  wire [7:0] rom__T_729_addr;
  wire  rom__T_729_mask;
  wire  rom__T_729_en;
  wire [7:0] rom__T_732_data;
  wire [7:0] rom__T_732_addr;
  wire  rom__T_732_mask;
  wire  rom__T_732_en;
  wire [7:0] rom__T_736_data;
  wire [7:0] rom__T_736_addr;
  wire  rom__T_736_mask;
  wire  rom__T_736_en;
  wire [7:0] rom__T_739_data;
  wire [7:0] rom__T_739_addr;
  wire  rom__T_739_mask;
  wire  rom__T_739_en;
  wire [7:0] rom__T_742_data;
  wire [7:0] rom__T_742_addr;
  wire  rom__T_742_mask;
  wire  rom__T_742_en;
  wire [7:0] rom__T_745_data;
  wire [7:0] rom__T_745_addr;
  wire  rom__T_745_mask;
  wire  rom__T_745_en;
  wire [7:0] rom__T_749_data;
  wire [7:0] rom__T_749_addr;
  wire  rom__T_749_mask;
  wire  rom__T_749_en;
  wire [7:0] rom__T_752_data;
  wire [7:0] rom__T_752_addr;
  wire  rom__T_752_mask;
  wire  rom__T_752_en;
  wire [7:0] rom__T_755_data;
  wire [7:0] rom__T_755_addr;
  wire  rom__T_755_mask;
  wire  rom__T_755_en;
  wire [7:0] rom__T_758_data;
  wire [7:0] rom__T_758_addr;
  wire  rom__T_758_mask;
  wire  rom__T_758_en;
  wire [7:0] rom__T_762_data;
  wire [7:0] rom__T_762_addr;
  wire  rom__T_762_mask;
  wire  rom__T_762_en;
  wire [7:0] rom__T_765_data;
  wire [7:0] rom__T_765_addr;
  wire  rom__T_765_mask;
  wire  rom__T_765_en;
  wire [7:0] rom__T_768_data;
  wire [7:0] rom__T_768_addr;
  wire  rom__T_768_mask;
  wire  rom__T_768_en;
  wire [7:0] rom__T_771_data;
  wire [7:0] rom__T_771_addr;
  wire  rom__T_771_mask;
  wire  rom__T_771_en;
  wire [7:0] rom__T_775_data;
  wire [7:0] rom__T_775_addr;
  wire  rom__T_775_mask;
  wire  rom__T_775_en;
  wire [7:0] rom__T_778_data;
  wire [7:0] rom__T_778_addr;
  wire  rom__T_778_mask;
  wire  rom__T_778_en;
  wire [7:0] rom__T_781_data;
  wire [7:0] rom__T_781_addr;
  wire  rom__T_781_mask;
  wire  rom__T_781_en;
  wire [7:0] rom__T_784_data;
  wire [7:0] rom__T_784_addr;
  wire  rom__T_784_mask;
  wire  rom__T_784_en;
  wire [32:0] _T_787;
  wire [31:0] _T_788;
  wire [7:0] _T_789;
  wire [32:0] _T_792;
  wire [31:0] _T_793;
  wire [7:0] _T_794;
  wire [32:0] _T_797;
  wire [31:0] _T_798;
  wire [7:0] _T_799;
  wire [7:0] _T_801;
  wire [15:0] _T_803;
  wire [15:0] _T_804;
  wire [31:0] _T_805;
  assign io_inst = _T_805;
  assign rom__T_790_addr = _T_789;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rom__T_790_data = rom[rom__T_790_addr];
  `else
  assign rom__T_790_data = rom__T_790_addr >= 8'hf0 ? _GEN_1[7:0] : rom[rom__T_790_addr];
  `endif
  assign rom__T_795_addr = _T_794;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rom__T_795_data = rom[rom__T_795_addr];
  `else
  assign rom__T_795_data = rom__T_795_addr >= 8'hf0 ? _GEN_2[7:0] : rom[rom__T_795_addr];
  `endif
  assign rom__T_800_addr = _T_799;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rom__T_800_data = rom[rom__T_800_addr];
  `else
  assign rom__T_800_data = rom__T_800_addr >= 8'hf0 ? _GEN_3[7:0] : rom[rom__T_800_addr];
  `endif
  assign rom__T_802_addr = _T_801;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rom__T_802_data = rom[rom__T_802_addr];
  `else
  assign rom__T_802_data = rom__T_802_addr >= 8'hf0 ? _GEN_4[7:0] : rom[rom__T_802_addr];
  `endif
  assign rom__T_8_data = 8'h7f;
  assign rom__T_8_addr = 8'h0;
  assign rom__T_8_mask = 1'h1;
  assign rom__T_8_en = 1'h1;
  assign rom__T_11_data = 8'h45;
  assign rom__T_11_addr = 8'h1;
  assign rom__T_11_mask = 1'h1;
  assign rom__T_11_en = 1'h1;
  assign rom__T_14_data = 8'h4c;
  assign rom__T_14_addr = 8'h2;
  assign rom__T_14_mask = 1'h1;
  assign rom__T_14_en = 1'h1;
  assign rom__T_17_data = 8'h46;
  assign rom__T_17_addr = 8'h3;
  assign rom__T_17_mask = 1'h1;
  assign rom__T_17_en = 1'h1;
  assign rom__T_21_data = 8'h1;
  assign rom__T_21_addr = 8'h4;
  assign rom__T_21_mask = 1'h1;
  assign rom__T_21_en = 1'h1;
  assign rom__T_24_data = 8'h1;
  assign rom__T_24_addr = 8'h5;
  assign rom__T_24_mask = 1'h1;
  assign rom__T_24_en = 1'h1;
  assign rom__T_27_data = 8'h1;
  assign rom__T_27_addr = 8'h6;
  assign rom__T_27_mask = 1'h1;
  assign rom__T_27_en = 1'h1;
  assign rom__T_30_data = 8'h0;
  assign rom__T_30_addr = 8'h7;
  assign rom__T_30_mask = 1'h1;
  assign rom__T_30_en = 1'h1;
  assign rom__T_34_data = 8'h0;
  assign rom__T_34_addr = 8'h8;
  assign rom__T_34_mask = 1'h1;
  assign rom__T_34_en = 1'h1;
  assign rom__T_37_data = 8'h0;
  assign rom__T_37_addr = 8'h9;
  assign rom__T_37_mask = 1'h1;
  assign rom__T_37_en = 1'h1;
  assign rom__T_40_data = 8'h0;
  assign rom__T_40_addr = 8'ha;
  assign rom__T_40_mask = 1'h1;
  assign rom__T_40_en = 1'h1;
  assign rom__T_43_data = 8'h0;
  assign rom__T_43_addr = 8'hb;
  assign rom__T_43_mask = 1'h1;
  assign rom__T_43_en = 1'h1;
  assign rom__T_47_data = 8'h0;
  assign rom__T_47_addr = 8'hc;
  assign rom__T_47_mask = 1'h1;
  assign rom__T_47_en = 1'h1;
  assign rom__T_50_data = 8'h0;
  assign rom__T_50_addr = 8'hd;
  assign rom__T_50_mask = 1'h1;
  assign rom__T_50_en = 1'h1;
  assign rom__T_53_data = 8'h0;
  assign rom__T_53_addr = 8'he;
  assign rom__T_53_mask = 1'h1;
  assign rom__T_53_en = 1'h1;
  assign rom__T_56_data = 8'h0;
  assign rom__T_56_addr = 8'hf;
  assign rom__T_56_mask = 1'h1;
  assign rom__T_56_en = 1'h1;
  assign rom__T_60_data = 8'h2;
  assign rom__T_60_addr = 8'h10;
  assign rom__T_60_mask = 1'h1;
  assign rom__T_60_en = 1'h1;
  assign rom__T_63_data = 8'h0;
  assign rom__T_63_addr = 8'h11;
  assign rom__T_63_mask = 1'h1;
  assign rom__T_63_en = 1'h1;
  assign rom__T_66_data = 8'hf3;
  assign rom__T_66_addr = 8'h12;
  assign rom__T_66_mask = 1'h1;
  assign rom__T_66_en = 1'h1;
  assign rom__T_69_data = 8'h0;
  assign rom__T_69_addr = 8'h13;
  assign rom__T_69_mask = 1'h1;
  assign rom__T_69_en = 1'h1;
  assign rom__T_73_data = 8'h1;
  assign rom__T_73_addr = 8'h14;
  assign rom__T_73_mask = 1'h1;
  assign rom__T_73_en = 1'h1;
  assign rom__T_76_data = 8'h0;
  assign rom__T_76_addr = 8'h15;
  assign rom__T_76_mask = 1'h1;
  assign rom__T_76_en = 1'h1;
  assign rom__T_79_data = 8'h0;
  assign rom__T_79_addr = 8'h16;
  assign rom__T_79_mask = 1'h1;
  assign rom__T_79_en = 1'h1;
  assign rom__T_82_data = 8'h0;
  assign rom__T_82_addr = 8'h17;
  assign rom__T_82_mask = 1'h1;
  assign rom__T_82_en = 1'h1;
  assign rom__T_86_data = 8'h54;
  assign rom__T_86_addr = 8'h18;
  assign rom__T_86_mask = 1'h1;
  assign rom__T_86_en = 1'h1;
  assign rom__T_89_data = 8'h0;
  assign rom__T_89_addr = 8'h19;
  assign rom__T_89_mask = 1'h1;
  assign rom__T_89_en = 1'h1;
  assign rom__T_92_data = 8'h1;
  assign rom__T_92_addr = 8'h1a;
  assign rom__T_92_mask = 1'h1;
  assign rom__T_92_en = 1'h1;
  assign rom__T_95_data = 8'h0;
  assign rom__T_95_addr = 8'h1b;
  assign rom__T_95_mask = 1'h1;
  assign rom__T_95_en = 1'h1;
  assign rom__T_99_data = 8'h34;
  assign rom__T_99_addr = 8'h1c;
  assign rom__T_99_mask = 1'h1;
  assign rom__T_99_en = 1'h1;
  assign rom__T_102_data = 8'h0;
  assign rom__T_102_addr = 8'h1d;
  assign rom__T_102_mask = 1'h1;
  assign rom__T_102_en = 1'h1;
  assign rom__T_105_data = 8'h0;
  assign rom__T_105_addr = 8'h1e;
  assign rom__T_105_mask = 1'h1;
  assign rom__T_105_en = 1'h1;
  assign rom__T_108_data = 8'h0;
  assign rom__T_108_addr = 8'h1f;
  assign rom__T_108_mask = 1'h1;
  assign rom__T_108_en = 1'h1;
  assign rom__T_112_data = 8'hdc;
  assign rom__T_112_addr = 8'h20;
  assign rom__T_112_mask = 1'h1;
  assign rom__T_112_en = 1'h1;
  assign rom__T_115_data = 8'h1;
  assign rom__T_115_addr = 8'h21;
  assign rom__T_115_mask = 1'h1;
  assign rom__T_115_en = 1'h1;
  assign rom__T_118_data = 8'h0;
  assign rom__T_118_addr = 8'h22;
  assign rom__T_118_mask = 1'h1;
  assign rom__T_118_en = 1'h1;
  assign rom__T_121_data = 8'h0;
  assign rom__T_121_addr = 8'h23;
  assign rom__T_121_mask = 1'h1;
  assign rom__T_121_en = 1'h1;
  assign rom__T_125_data = 8'h0;
  assign rom__T_125_addr = 8'h24;
  assign rom__T_125_mask = 1'h1;
  assign rom__T_125_en = 1'h1;
  assign rom__T_128_data = 8'h0;
  assign rom__T_128_addr = 8'h25;
  assign rom__T_128_mask = 1'h1;
  assign rom__T_128_en = 1'h1;
  assign rom__T_131_data = 8'h0;
  assign rom__T_131_addr = 8'h26;
  assign rom__T_131_mask = 1'h1;
  assign rom__T_131_en = 1'h1;
  assign rom__T_134_data = 8'h0;
  assign rom__T_134_addr = 8'h27;
  assign rom__T_134_mask = 1'h1;
  assign rom__T_134_en = 1'h1;
  assign rom__T_138_data = 8'h34;
  assign rom__T_138_addr = 8'h28;
  assign rom__T_138_mask = 1'h1;
  assign rom__T_138_en = 1'h1;
  assign rom__T_141_data = 8'h0;
  assign rom__T_141_addr = 8'h29;
  assign rom__T_141_mask = 1'h1;
  assign rom__T_141_en = 1'h1;
  assign rom__T_144_data = 8'h20;
  assign rom__T_144_addr = 8'h2a;
  assign rom__T_144_mask = 1'h1;
  assign rom__T_144_en = 1'h1;
  assign rom__T_147_data = 8'h0;
  assign rom__T_147_addr = 8'h2b;
  assign rom__T_147_mask = 1'h1;
  assign rom__T_147_en = 1'h1;
  assign rom__T_151_data = 8'h1;
  assign rom__T_151_addr = 8'h2c;
  assign rom__T_151_mask = 1'h1;
  assign rom__T_151_en = 1'h1;
  assign rom__T_154_data = 8'h0;
  assign rom__T_154_addr = 8'h2d;
  assign rom__T_154_mask = 1'h1;
  assign rom__T_154_en = 1'h1;
  assign rom__T_157_data = 8'h28;
  assign rom__T_157_addr = 8'h2e;
  assign rom__T_157_mask = 1'h1;
  assign rom__T_157_en = 1'h1;
  assign rom__T_160_data = 8'h0;
  assign rom__T_160_addr = 8'h2f;
  assign rom__T_160_mask = 1'h1;
  assign rom__T_160_en = 1'h1;
  assign rom__T_164_data = 8'h6;
  assign rom__T_164_addr = 8'h30;
  assign rom__T_164_mask = 1'h1;
  assign rom__T_164_en = 1'h1;
  assign rom__T_167_data = 8'h0;
  assign rom__T_167_addr = 8'h31;
  assign rom__T_167_mask = 1'h1;
  assign rom__T_167_en = 1'h1;
  assign rom__T_170_data = 8'h5;
  assign rom__T_170_addr = 8'h32;
  assign rom__T_170_mask = 1'h1;
  assign rom__T_170_en = 1'h1;
  assign rom__T_173_data = 8'h0;
  assign rom__T_173_addr = 8'h33;
  assign rom__T_173_mask = 1'h1;
  assign rom__T_173_en = 1'h1;
  assign rom__T_177_data = 8'h1;
  assign rom__T_177_addr = 8'h34;
  assign rom__T_177_mask = 1'h1;
  assign rom__T_177_en = 1'h1;
  assign rom__T_180_data = 8'h0;
  assign rom__T_180_addr = 8'h35;
  assign rom__T_180_mask = 1'h1;
  assign rom__T_180_en = 1'h1;
  assign rom__T_183_data = 8'h0;
  assign rom__T_183_addr = 8'h36;
  assign rom__T_183_mask = 1'h1;
  assign rom__T_183_en = 1'h1;
  assign rom__T_186_data = 8'h0;
  assign rom__T_186_addr = 8'h37;
  assign rom__T_186_mask = 1'h1;
  assign rom__T_186_en = 1'h1;
  assign rom__T_190_data = 8'h0;
  assign rom__T_190_addr = 8'h38;
  assign rom__T_190_mask = 1'h1;
  assign rom__T_190_en = 1'h1;
  assign rom__T_193_data = 8'h0;
  assign rom__T_193_addr = 8'h39;
  assign rom__T_193_mask = 1'h1;
  assign rom__T_193_en = 1'h1;
  assign rom__T_196_data = 8'h0;
  assign rom__T_196_addr = 8'h3a;
  assign rom__T_196_mask = 1'h1;
  assign rom__T_196_en = 1'h1;
  assign rom__T_199_data = 8'h0;
  assign rom__T_199_addr = 8'h3b;
  assign rom__T_199_mask = 1'h1;
  assign rom__T_199_en = 1'h1;
  assign rom__T_203_data = 8'h0;
  assign rom__T_203_addr = 8'h3c;
  assign rom__T_203_mask = 1'h1;
  assign rom__T_203_en = 1'h1;
  assign rom__T_206_data = 8'h0;
  assign rom__T_206_addr = 8'h3d;
  assign rom__T_206_mask = 1'h1;
  assign rom__T_206_en = 1'h1;
  assign rom__T_209_data = 8'h1;
  assign rom__T_209_addr = 8'h3e;
  assign rom__T_209_mask = 1'h1;
  assign rom__T_209_en = 1'h1;
  assign rom__T_212_data = 8'h0;
  assign rom__T_212_addr = 8'h3f;
  assign rom__T_212_mask = 1'h1;
  assign rom__T_212_en = 1'h1;
  assign rom__T_216_data = 8'h0;
  assign rom__T_216_addr = 8'h40;
  assign rom__T_216_mask = 1'h1;
  assign rom__T_216_en = 1'h1;
  assign rom__T_219_data = 8'h0;
  assign rom__T_219_addr = 8'h41;
  assign rom__T_219_mask = 1'h1;
  assign rom__T_219_en = 1'h1;
  assign rom__T_222_data = 8'h1;
  assign rom__T_222_addr = 8'h42;
  assign rom__T_222_mask = 1'h1;
  assign rom__T_222_en = 1'h1;
  assign rom__T_225_data = 8'h0;
  assign rom__T_225_addr = 8'h43;
  assign rom__T_225_mask = 1'h1;
  assign rom__T_225_en = 1'h1;
  assign rom__T_229_data = 8'hcc;
  assign rom__T_229_addr = 8'h44;
  assign rom__T_229_mask = 1'h1;
  assign rom__T_229_en = 1'h1;
  assign rom__T_232_data = 8'h0;
  assign rom__T_232_addr = 8'h45;
  assign rom__T_232_mask = 1'h1;
  assign rom__T_232_en = 1'h1;
  assign rom__T_235_data = 8'h0;
  assign rom__T_235_addr = 8'h46;
  assign rom__T_235_mask = 1'h1;
  assign rom__T_235_en = 1'h1;
  assign rom__T_238_data = 8'h0;
  assign rom__T_238_addr = 8'h47;
  assign rom__T_238_mask = 1'h1;
  assign rom__T_238_en = 1'h1;
  assign rom__T_242_data = 8'hcc;
  assign rom__T_242_addr = 8'h48;
  assign rom__T_242_mask = 1'h1;
  assign rom__T_242_en = 1'h1;
  assign rom__T_245_data = 8'h0;
  assign rom__T_245_addr = 8'h49;
  assign rom__T_245_mask = 1'h1;
  assign rom__T_245_en = 1'h1;
  assign rom__T_248_data = 8'h0;
  assign rom__T_248_addr = 8'h4a;
  assign rom__T_248_mask = 1'h1;
  assign rom__T_248_en = 1'h1;
  assign rom__T_251_data = 8'h0;
  assign rom__T_251_addr = 8'h4b;
  assign rom__T_251_mask = 1'h1;
  assign rom__T_251_en = 1'h1;
  assign rom__T_255_data = 8'h5;
  assign rom__T_255_addr = 8'h4c;
  assign rom__T_255_mask = 1'h1;
  assign rom__T_255_en = 1'h1;
  assign rom__T_258_data = 8'h0;
  assign rom__T_258_addr = 8'h4d;
  assign rom__T_258_mask = 1'h1;
  assign rom__T_258_en = 1'h1;
  assign rom__T_261_data = 8'h0;
  assign rom__T_261_addr = 8'h4e;
  assign rom__T_261_mask = 1'h1;
  assign rom__T_261_en = 1'h1;
  assign rom__T_264_data = 8'h0;
  assign rom__T_264_addr = 8'h4f;
  assign rom__T_264_mask = 1'h1;
  assign rom__T_264_en = 1'h1;
  assign rom__T_268_data = 8'h0;
  assign rom__T_268_addr = 8'h50;
  assign rom__T_268_mask = 1'h1;
  assign rom__T_268_en = 1'h1;
  assign rom__T_271_data = 8'h10;
  assign rom__T_271_addr = 8'h51;
  assign rom__T_271_mask = 1'h1;
  assign rom__T_271_en = 1'h1;
  assign rom__T_274_data = 8'h0;
  assign rom__T_274_addr = 8'h52;
  assign rom__T_274_mask = 1'h1;
  assign rom__T_274_en = 1'h1;
  assign rom__T_277_data = 8'h0;
  assign rom__T_277_addr = 8'h53;
  assign rom__T_277_mask = 1'h1;
  assign rom__T_277_en = 1'h1;
  assign rom__T_281_data = 8'h13;
  assign rom__T_281_addr = 8'h54;
  assign rom__T_281_mask = 1'h1;
  assign rom__T_281_en = 1'h1;
  assign rom__T_284_data = 8'h3;
  assign rom__T_284_addr = 8'h55;
  assign rom__T_284_mask = 1'h1;
  assign rom__T_284_en = 1'h1;
  assign rom__T_287_data = 8'h10;
  assign rom__T_287_addr = 8'h56;
  assign rom__T_287_mask = 1'h1;
  assign rom__T_287_en = 1'h1;
  assign rom__T_290_data = 8'h40;
  assign rom__T_290_addr = 8'h57;
  assign rom__T_290_mask = 1'h1;
  assign rom__T_290_en = 1'h1;
  assign rom__T_294_data = 8'h93;
  assign rom__T_294_addr = 8'h58;
  assign rom__T_294_mask = 1'h1;
  assign rom__T_294_en = 1'h1;
  assign rom__T_297_data = 8'h2;
  assign rom__T_297_addr = 8'h59;
  assign rom__T_297_mask = 1'h1;
  assign rom__T_297_en = 1'h1;
  assign rom__T_300_data = 8'h80;
  assign rom__T_300_addr = 8'h5a;
  assign rom__T_300_mask = 1'h1;
  assign rom__T_300_en = 1'h1;
  assign rom__T_303_data = 8'h6;
  assign rom__T_303_addr = 8'h5b;
  assign rom__T_303_mask = 1'h1;
  assign rom__T_303_en = 1'h1;
  assign rom__T_307_data = 8'h23;
  assign rom__T_307_addr = 8'h5c;
  assign rom__T_307_mask = 1'h1;
  assign rom__T_307_en = 1'h1;
  assign rom__T_310_data = 8'h20;
  assign rom__T_310_addr = 8'h5d;
  assign rom__T_310_mask = 1'h1;
  assign rom__T_310_en = 1'h1;
  assign rom__T_313_data = 8'h53;
  assign rom__T_313_addr = 8'h5e;
  assign rom__T_313_mask = 1'h1;
  assign rom__T_313_en = 1'h1;
  assign rom__T_316_data = 8'h0;
  assign rom__T_316_addr = 8'h5f;
  assign rom__T_316_mask = 1'h1;
  assign rom__T_316_en = 1'h1;
  assign rom__T_320_data = 8'h93;
  assign rom__T_320_addr = 8'h60;
  assign rom__T_320_mask = 1'h1;
  assign rom__T_320_en = 1'h1;
  assign rom__T_323_data = 8'h2;
  assign rom__T_323_addr = 8'h61;
  assign rom__T_323_mask = 1'h1;
  assign rom__T_323_en = 1'h1;
  assign rom__T_326_data = 8'h50;
  assign rom__T_326_addr = 8'h62;
  assign rom__T_326_mask = 1'h1;
  assign rom__T_326_en = 1'h1;
  assign rom__T_329_data = 8'h6;
  assign rom__T_329_addr = 8'h63;
  assign rom__T_329_mask = 1'h1;
  assign rom__T_329_en = 1'h1;
  assign rom__T_333_data = 8'h23;
  assign rom__T_333_addr = 8'h64;
  assign rom__T_333_mask = 1'h1;
  assign rom__T_333_en = 1'h1;
  assign rom__T_336_data = 8'h20;
  assign rom__T_336_addr = 8'h65;
  assign rom__T_336_mask = 1'h1;
  assign rom__T_336_en = 1'h1;
  assign rom__T_339_data = 8'h53;
  assign rom__T_339_addr = 8'h66;
  assign rom__T_339_mask = 1'h1;
  assign rom__T_339_en = 1'h1;
  assign rom__T_342_data = 8'h0;
  assign rom__T_342_addr = 8'h67;
  assign rom__T_342_mask = 1'h1;
  assign rom__T_342_en = 1'h1;
  assign rom__T_346_data = 8'h93;
  assign rom__T_346_addr = 8'h68;
  assign rom__T_346_mask = 1'h1;
  assign rom__T_346_en = 1'h1;
  assign rom__T_349_data = 8'h2;
  assign rom__T_349_addr = 8'h69;
  assign rom__T_349_mask = 1'h1;
  assign rom__T_349_en = 1'h1;
  assign rom__T_352_data = 8'hc0;
  assign rom__T_352_addr = 8'h6a;
  assign rom__T_352_mask = 1'h1;
  assign rom__T_352_en = 1'h1;
  assign rom__T_355_data = 8'h6;
  assign rom__T_355_addr = 8'h6b;
  assign rom__T_355_mask = 1'h1;
  assign rom__T_355_en = 1'h1;
  assign rom__T_359_data = 8'h23;
  assign rom__T_359_addr = 8'h6c;
  assign rom__T_359_mask = 1'h1;
  assign rom__T_359_en = 1'h1;
  assign rom__T_362_data = 8'h20;
  assign rom__T_362_addr = 8'h6d;
  assign rom__T_362_mask = 1'h1;
  assign rom__T_362_en = 1'h1;
  assign rom__T_365_data = 8'h53;
  assign rom__T_365_addr = 8'h6e;
  assign rom__T_365_mask = 1'h1;
  assign rom__T_365_en = 1'h1;
  assign rom__T_368_data = 8'h0;
  assign rom__T_368_addr = 8'h6f;
  assign rom__T_368_mask = 1'h1;
  assign rom__T_368_en = 1'h1;
  assign rom__T_372_data = 8'h93;
  assign rom__T_372_addr = 8'h70;
  assign rom__T_372_mask = 1'h1;
  assign rom__T_372_en = 1'h1;
  assign rom__T_375_data = 8'h2;
  assign rom__T_375_addr = 8'h71;
  assign rom__T_375_mask = 1'h1;
  assign rom__T_375_en = 1'h1;
  assign rom__T_378_data = 8'hc0;
  assign rom__T_378_addr = 8'h72;
  assign rom__T_378_mask = 1'h1;
  assign rom__T_378_en = 1'h1;
  assign rom__T_381_data = 8'h6;
  assign rom__T_381_addr = 8'h73;
  assign rom__T_381_mask = 1'h1;
  assign rom__T_381_en = 1'h1;
  assign rom__T_385_data = 8'h23;
  assign rom__T_385_addr = 8'h74;
  assign rom__T_385_mask = 1'h1;
  assign rom__T_385_en = 1'h1;
  assign rom__T_388_data = 8'h20;
  assign rom__T_388_addr = 8'h75;
  assign rom__T_388_mask = 1'h1;
  assign rom__T_388_en = 1'h1;
  assign rom__T_391_data = 8'h53;
  assign rom__T_391_addr = 8'h76;
  assign rom__T_391_mask = 1'h1;
  assign rom__T_391_en = 1'h1;
  assign rom__T_394_data = 8'h0;
  assign rom__T_394_addr = 8'h77;
  assign rom__T_394_mask = 1'h1;
  assign rom__T_394_en = 1'h1;
  assign rom__T_398_data = 8'h93;
  assign rom__T_398_addr = 8'h78;
  assign rom__T_398_mask = 1'h1;
  assign rom__T_398_en = 1'h1;
  assign rom__T_401_data = 8'h2;
  assign rom__T_401_addr = 8'h79;
  assign rom__T_401_mask = 1'h1;
  assign rom__T_401_en = 1'h1;
  assign rom__T_404_data = 8'hf0;
  assign rom__T_404_addr = 8'h7a;
  assign rom__T_404_mask = 1'h1;
  assign rom__T_404_en = 1'h1;
  assign rom__T_407_data = 8'h6;
  assign rom__T_407_addr = 8'h7b;
  assign rom__T_407_mask = 1'h1;
  assign rom__T_407_en = 1'h1;
  assign rom__T_411_data = 8'h23;
  assign rom__T_411_addr = 8'h7c;
  assign rom__T_411_mask = 1'h1;
  assign rom__T_411_en = 1'h1;
  assign rom__T_414_data = 8'h20;
  assign rom__T_414_addr = 8'h7d;
  assign rom__T_414_mask = 1'h1;
  assign rom__T_414_en = 1'h1;
  assign rom__T_417_data = 8'h53;
  assign rom__T_417_addr = 8'h7e;
  assign rom__T_417_mask = 1'h1;
  assign rom__T_417_en = 1'h1;
  assign rom__T_420_data = 8'h0;
  assign rom__T_420_addr = 8'h7f;
  assign rom__T_420_mask = 1'h1;
  assign rom__T_420_en = 1'h1;
  assign rom__T_424_data = 8'h93;
  assign rom__T_424_addr = 8'h80;
  assign rom__T_424_mask = 1'h1;
  assign rom__T_424_en = 1'h1;
  assign rom__T_427_data = 8'h2;
  assign rom__T_427_addr = 8'h81;
  assign rom__T_427_mask = 1'h1;
  assign rom__T_427_en = 1'h1;
  assign rom__T_430_data = 8'h0;
  assign rom__T_430_addr = 8'h82;
  assign rom__T_430_mask = 1'h1;
  assign rom__T_430_en = 1'h1;
  assign rom__T_433_data = 8'h2;
  assign rom__T_433_addr = 8'h83;
  assign rom__T_433_mask = 1'h1;
  assign rom__T_433_en = 1'h1;
  assign rom__T_437_data = 8'h23;
  assign rom__T_437_addr = 8'h84;
  assign rom__T_437_mask = 1'h1;
  assign rom__T_437_en = 1'h1;
  assign rom__T_440_data = 8'h20;
  assign rom__T_440_addr = 8'h85;
  assign rom__T_440_mask = 1'h1;
  assign rom__T_440_en = 1'h1;
  assign rom__T_443_data = 8'h53;
  assign rom__T_443_addr = 8'h86;
  assign rom__T_443_mask = 1'h1;
  assign rom__T_443_en = 1'h1;
  assign rom__T_446_data = 8'h0;
  assign rom__T_446_addr = 8'h87;
  assign rom__T_446_mask = 1'h1;
  assign rom__T_446_en = 1'h1;
  assign rom__T_450_data = 8'h93;
  assign rom__T_450_addr = 8'h88;
  assign rom__T_450_mask = 1'h1;
  assign rom__T_450_en = 1'h1;
  assign rom__T_453_data = 8'h2;
  assign rom__T_453_addr = 8'h89;
  assign rom__T_453_mask = 1'h1;
  assign rom__T_453_en = 1'h1;
  assign rom__T_456_data = 8'h70;
  assign rom__T_456_addr = 8'h8a;
  assign rom__T_456_mask = 1'h1;
  assign rom__T_456_en = 1'h1;
  assign rom__T_459_data = 8'h7;
  assign rom__T_459_addr = 8'h8b;
  assign rom__T_459_mask = 1'h1;
  assign rom__T_459_en = 1'h1;
  assign rom__T_463_data = 8'h23;
  assign rom__T_463_addr = 8'h8c;
  assign rom__T_463_mask = 1'h1;
  assign rom__T_463_en = 1'h1;
  assign rom__T_466_data = 8'h20;
  assign rom__T_466_addr = 8'h8d;
  assign rom__T_466_mask = 1'h1;
  assign rom__T_466_en = 1'h1;
  assign rom__T_469_data = 8'h53;
  assign rom__T_469_addr = 8'h8e;
  assign rom__T_469_mask = 1'h1;
  assign rom__T_469_en = 1'h1;
  assign rom__T_472_data = 8'h0;
  assign rom__T_472_addr = 8'h8f;
  assign rom__T_472_mask = 1'h1;
  assign rom__T_472_en = 1'h1;
  assign rom__T_476_data = 8'h93;
  assign rom__T_476_addr = 8'h90;
  assign rom__T_476_mask = 1'h1;
  assign rom__T_476_en = 1'h1;
  assign rom__T_479_data = 8'h2;
  assign rom__T_479_addr = 8'h91;
  assign rom__T_479_mask = 1'h1;
  assign rom__T_479_en = 1'h1;
  assign rom__T_482_data = 8'hf0;
  assign rom__T_482_addr = 8'h92;
  assign rom__T_482_mask = 1'h1;
  assign rom__T_482_en = 1'h1;
  assign rom__T_485_data = 8'h6;
  assign rom__T_485_addr = 8'h93;
  assign rom__T_485_mask = 1'h1;
  assign rom__T_485_en = 1'h1;
  assign rom__T_489_data = 8'h23;
  assign rom__T_489_addr = 8'h94;
  assign rom__T_489_mask = 1'h1;
  assign rom__T_489_en = 1'h1;
  assign rom__T_492_data = 8'h20;
  assign rom__T_492_addr = 8'h95;
  assign rom__T_492_mask = 1'h1;
  assign rom__T_492_en = 1'h1;
  assign rom__T_495_data = 8'h53;
  assign rom__T_495_addr = 8'h96;
  assign rom__T_495_mask = 1'h1;
  assign rom__T_495_en = 1'h1;
  assign rom__T_498_data = 8'h0;
  assign rom__T_498_addr = 8'h97;
  assign rom__T_498_mask = 1'h1;
  assign rom__T_498_en = 1'h1;
  assign rom__T_502_data = 8'h93;
  assign rom__T_502_addr = 8'h98;
  assign rom__T_502_mask = 1'h1;
  assign rom__T_502_en = 1'h1;
  assign rom__T_505_data = 8'h2;
  assign rom__T_505_addr = 8'h99;
  assign rom__T_505_mask = 1'h1;
  assign rom__T_505_en = 1'h1;
  assign rom__T_508_data = 8'h20;
  assign rom__T_508_addr = 8'h9a;
  assign rom__T_508_mask = 1'h1;
  assign rom__T_508_en = 1'h1;
  assign rom__T_511_data = 8'h7;
  assign rom__T_511_addr = 8'h9b;
  assign rom__T_511_mask = 1'h1;
  assign rom__T_511_en = 1'h1;
  assign rom__T_515_data = 8'h23;
  assign rom__T_515_addr = 8'h9c;
  assign rom__T_515_mask = 1'h1;
  assign rom__T_515_en = 1'h1;
  assign rom__T_518_data = 8'h20;
  assign rom__T_518_addr = 8'h9d;
  assign rom__T_518_mask = 1'h1;
  assign rom__T_518_en = 1'h1;
  assign rom__T_521_data = 8'h53;
  assign rom__T_521_addr = 8'h9e;
  assign rom__T_521_mask = 1'h1;
  assign rom__T_521_en = 1'h1;
  assign rom__T_524_data = 8'h0;
  assign rom__T_524_addr = 8'h9f;
  assign rom__T_524_mask = 1'h1;
  assign rom__T_524_en = 1'h1;
  assign rom__T_528_data = 8'h93;
  assign rom__T_528_addr = 8'ha0;
  assign rom__T_528_mask = 1'h1;
  assign rom__T_528_en = 1'h1;
  assign rom__T_531_data = 8'h2;
  assign rom__T_531_addr = 8'ha1;
  assign rom__T_531_mask = 1'h1;
  assign rom__T_531_en = 1'h1;
  assign rom__T_534_data = 8'hc0;
  assign rom__T_534_addr = 8'ha2;
  assign rom__T_534_mask = 1'h1;
  assign rom__T_534_en = 1'h1;
  assign rom__T_537_data = 8'h6;
  assign rom__T_537_addr = 8'ha3;
  assign rom__T_537_mask = 1'h1;
  assign rom__T_537_en = 1'h1;
  assign rom__T_541_data = 8'h23;
  assign rom__T_541_addr = 8'ha4;
  assign rom__T_541_mask = 1'h1;
  assign rom__T_541_en = 1'h1;
  assign rom__T_544_data = 8'h20;
  assign rom__T_544_addr = 8'ha5;
  assign rom__T_544_mask = 1'h1;
  assign rom__T_544_en = 1'h1;
  assign rom__T_547_data = 8'h53;
  assign rom__T_547_addr = 8'ha6;
  assign rom__T_547_mask = 1'h1;
  assign rom__T_547_en = 1'h1;
  assign rom__T_550_data = 8'h0;
  assign rom__T_550_addr = 8'ha7;
  assign rom__T_550_mask = 1'h1;
  assign rom__T_550_en = 1'h1;
  assign rom__T_554_data = 8'h93;
  assign rom__T_554_addr = 8'ha8;
  assign rom__T_554_mask = 1'h1;
  assign rom__T_554_en = 1'h1;
  assign rom__T_557_data = 8'h2;
  assign rom__T_557_addr = 8'ha9;
  assign rom__T_557_mask = 1'h1;
  assign rom__T_557_en = 1'h1;
  assign rom__T_560_data = 8'h40;
  assign rom__T_560_addr = 8'haa;
  assign rom__T_560_mask = 1'h1;
  assign rom__T_560_en = 1'h1;
  assign rom__T_563_data = 8'h6;
  assign rom__T_563_addr = 8'hab;
  assign rom__T_563_mask = 1'h1;
  assign rom__T_563_en = 1'h1;
  assign rom__T_567_data = 8'h23;
  assign rom__T_567_addr = 8'hac;
  assign rom__T_567_mask = 1'h1;
  assign rom__T_567_en = 1'h1;
  assign rom__T_570_data = 8'h20;
  assign rom__T_570_addr = 8'had;
  assign rom__T_570_mask = 1'h1;
  assign rom__T_570_en = 1'h1;
  assign rom__T_573_data = 8'h53;
  assign rom__T_573_addr = 8'hae;
  assign rom__T_573_mask = 1'h1;
  assign rom__T_573_en = 1'h1;
  assign rom__T_576_data = 8'h0;
  assign rom__T_576_addr = 8'haf;
  assign rom__T_576_mask = 1'h1;
  assign rom__T_576_en = 1'h1;
  assign rom__T_580_data = 8'h93;
  assign rom__T_580_addr = 8'hb0;
  assign rom__T_580_mask = 1'h1;
  assign rom__T_580_en = 1'h1;
  assign rom__T_583_data = 8'h2;
  assign rom__T_583_addr = 8'hb1;
  assign rom__T_583_mask = 1'h1;
  assign rom__T_583_en = 1'h1;
  assign rom__T_586_data = 8'h10;
  assign rom__T_586_addr = 8'hb2;
  assign rom__T_586_mask = 1'h1;
  assign rom__T_586_en = 1'h1;
  assign rom__T_589_data = 8'h2;
  assign rom__T_589_addr = 8'hb3;
  assign rom__T_589_mask = 1'h1;
  assign rom__T_589_en = 1'h1;
  assign rom__T_593_data = 8'h23;
  assign rom__T_593_addr = 8'hb4;
  assign rom__T_593_mask = 1'h1;
  assign rom__T_593_en = 1'h1;
  assign rom__T_596_data = 8'h20;
  assign rom__T_596_addr = 8'hb5;
  assign rom__T_596_mask = 1'h1;
  assign rom__T_596_en = 1'h1;
  assign rom__T_599_data = 8'h53;
  assign rom__T_599_addr = 8'hb6;
  assign rom__T_599_mask = 1'h1;
  assign rom__T_599_en = 1'h1;
  assign rom__T_602_data = 8'h0;
  assign rom__T_602_addr = 8'hb7;
  assign rom__T_602_mask = 1'h1;
  assign rom__T_602_en = 1'h1;
  assign rom__T_606_data = 8'h93;
  assign rom__T_606_addr = 8'hb8;
  assign rom__T_606_mask = 1'h1;
  assign rom__T_606_en = 1'h1;
  assign rom__T_609_data = 8'h2;
  assign rom__T_609_addr = 8'hb9;
  assign rom__T_609_mask = 1'h1;
  assign rom__T_609_en = 1'h1;
  assign rom__T_612_data = 8'ha0;
  assign rom__T_612_addr = 8'hba;
  assign rom__T_612_mask = 1'h1;
  assign rom__T_612_en = 1'h1;
  assign rom__T_615_data = 8'h0;
  assign rom__T_615_addr = 8'hbb;
  assign rom__T_615_mask = 1'h1;
  assign rom__T_615_en = 1'h1;
  assign rom__T_619_data = 8'h23;
  assign rom__T_619_addr = 8'hbc;
  assign rom__T_619_mask = 1'h1;
  assign rom__T_619_en = 1'h1;
  assign rom__T_622_data = 8'h20;
  assign rom__T_622_addr = 8'hbd;
  assign rom__T_622_mask = 1'h1;
  assign rom__T_622_en = 1'h1;
  assign rom__T_625_data = 8'h53;
  assign rom__T_625_addr = 8'hbe;
  assign rom__T_625_mask = 1'h1;
  assign rom__T_625_en = 1'h1;
  assign rom__T_628_data = 8'h0;
  assign rom__T_628_addr = 8'hbf;
  assign rom__T_628_mask = 1'h1;
  assign rom__T_628_en = 1'h1;
  assign rom__T_632_data = 8'h93;
  assign rom__T_632_addr = 8'hc0;
  assign rom__T_632_mask = 1'h1;
  assign rom__T_632_en = 1'h1;
  assign rom__T_635_data = 8'h2;
  assign rom__T_635_addr = 8'hc1;
  assign rom__T_635_mask = 1'h1;
  assign rom__T_635_en = 1'h1;
  assign rom__T_638_data = 8'hd0;
  assign rom__T_638_addr = 8'hc2;
  assign rom__T_638_mask = 1'h1;
  assign rom__T_638_en = 1'h1;
  assign rom__T_641_data = 8'h0;
  assign rom__T_641_addr = 8'hc3;
  assign rom__T_641_mask = 1'h1;
  assign rom__T_641_en = 1'h1;
  assign rom__T_645_data = 8'h23;
  assign rom__T_645_addr = 8'hc4;
  assign rom__T_645_mask = 1'h1;
  assign rom__T_645_en = 1'h1;
  assign rom__T_648_data = 8'h20;
  assign rom__T_648_addr = 8'hc5;
  assign rom__T_648_mask = 1'h1;
  assign rom__T_648_en = 1'h1;
  assign rom__T_651_data = 8'h53;
  assign rom__T_651_addr = 8'hc6;
  assign rom__T_651_mask = 1'h1;
  assign rom__T_651_en = 1'h1;
  assign rom__T_654_data = 8'h0;
  assign rom__T_654_addr = 8'hc7;
  assign rom__T_654_mask = 1'h1;
  assign rom__T_654_en = 1'h1;
  assign rom__T_658_data = 8'h67;
  assign rom__T_658_addr = 8'hc8;
  assign rom__T_658_mask = 1'h1;
  assign rom__T_658_en = 1'h1;
  assign rom__T_661_data = 8'h80;
  assign rom__T_661_addr = 8'hc9;
  assign rom__T_661_mask = 1'h1;
  assign rom__T_661_en = 1'h1;
  assign rom__T_664_data = 8'h0;
  assign rom__T_664_addr = 8'hca;
  assign rom__T_664_mask = 1'h1;
  assign rom__T_664_en = 1'h1;
  assign rom__T_667_data = 8'h0;
  assign rom__T_667_addr = 8'hcb;
  assign rom__T_667_mask = 1'h1;
  assign rom__T_667_en = 1'h1;
  assign rom__T_671_data = 8'h0;
  assign rom__T_671_addr = 8'hcc;
  assign rom__T_671_mask = 1'h1;
  assign rom__T_671_en = 1'h1;
  assign rom__T_674_data = 8'h0;
  assign rom__T_674_addr = 8'hcd;
  assign rom__T_674_mask = 1'h1;
  assign rom__T_674_en = 1'h1;
  assign rom__T_677_data = 8'h0;
  assign rom__T_677_addr = 8'hce;
  assign rom__T_677_mask = 1'h1;
  assign rom__T_677_en = 1'h1;
  assign rom__T_680_data = 8'h0;
  assign rom__T_680_addr = 8'hcf;
  assign rom__T_680_mask = 1'h1;
  assign rom__T_680_en = 1'h1;
  assign rom__T_684_data = 8'h0;
  assign rom__T_684_addr = 8'hd0;
  assign rom__T_684_mask = 1'h1;
  assign rom__T_684_en = 1'h1;
  assign rom__T_687_data = 8'h0;
  assign rom__T_687_addr = 8'hd1;
  assign rom__T_687_mask = 1'h1;
  assign rom__T_687_en = 1'h1;
  assign rom__T_690_data = 8'h0;
  assign rom__T_690_addr = 8'hd2;
  assign rom__T_690_mask = 1'h1;
  assign rom__T_690_en = 1'h1;
  assign rom__T_693_data = 8'h0;
  assign rom__T_693_addr = 8'hd3;
  assign rom__T_693_mask = 1'h1;
  assign rom__T_693_en = 1'h1;
  assign rom__T_697_data = 8'h0;
  assign rom__T_697_addr = 8'hd4;
  assign rom__T_697_mask = 1'h1;
  assign rom__T_697_en = 1'h1;
  assign rom__T_700_data = 8'h0;
  assign rom__T_700_addr = 8'hd5;
  assign rom__T_700_mask = 1'h1;
  assign rom__T_700_en = 1'h1;
  assign rom__T_703_data = 8'h0;
  assign rom__T_703_addr = 8'hd6;
  assign rom__T_703_mask = 1'h1;
  assign rom__T_703_en = 1'h1;
  assign rom__T_706_data = 8'h0;
  assign rom__T_706_addr = 8'hd7;
  assign rom__T_706_mask = 1'h1;
  assign rom__T_706_en = 1'h1;
  assign rom__T_710_data = 8'h0;
  assign rom__T_710_addr = 8'hd8;
  assign rom__T_710_mask = 1'h1;
  assign rom__T_710_en = 1'h1;
  assign rom__T_713_data = 8'h0;
  assign rom__T_713_addr = 8'hd9;
  assign rom__T_713_mask = 1'h1;
  assign rom__T_713_en = 1'h1;
  assign rom__T_716_data = 8'h0;
  assign rom__T_716_addr = 8'hda;
  assign rom__T_716_mask = 1'h1;
  assign rom__T_716_en = 1'h1;
  assign rom__T_719_data = 8'h0;
  assign rom__T_719_addr = 8'hdb;
  assign rom__T_719_mask = 1'h1;
  assign rom__T_719_en = 1'h1;
  assign rom__T_723_data = 8'h0;
  assign rom__T_723_addr = 8'hdc;
  assign rom__T_723_mask = 1'h1;
  assign rom__T_723_en = 1'h1;
  assign rom__T_726_data = 8'h0;
  assign rom__T_726_addr = 8'hdd;
  assign rom__T_726_mask = 1'h1;
  assign rom__T_726_en = 1'h1;
  assign rom__T_729_data = 8'h0;
  assign rom__T_729_addr = 8'hde;
  assign rom__T_729_mask = 1'h1;
  assign rom__T_729_en = 1'h1;
  assign rom__T_732_data = 8'h0;
  assign rom__T_732_addr = 8'hdf;
  assign rom__T_732_mask = 1'h1;
  assign rom__T_732_en = 1'h1;
  assign rom__T_736_data = 8'h0;
  assign rom__T_736_addr = 8'he0;
  assign rom__T_736_mask = 1'h1;
  assign rom__T_736_en = 1'h1;
  assign rom__T_739_data = 8'h0;
  assign rom__T_739_addr = 8'he1;
  assign rom__T_739_mask = 1'h1;
  assign rom__T_739_en = 1'h1;
  assign rom__T_742_data = 8'h0;
  assign rom__T_742_addr = 8'he2;
  assign rom__T_742_mask = 1'h1;
  assign rom__T_742_en = 1'h1;
  assign rom__T_745_data = 8'h0;
  assign rom__T_745_addr = 8'he3;
  assign rom__T_745_mask = 1'h1;
  assign rom__T_745_en = 1'h1;
  assign rom__T_749_data = 8'h0;
  assign rom__T_749_addr = 8'he4;
  assign rom__T_749_mask = 1'h1;
  assign rom__T_749_en = 1'h1;
  assign rom__T_752_data = 8'h0;
  assign rom__T_752_addr = 8'he5;
  assign rom__T_752_mask = 1'h1;
  assign rom__T_752_en = 1'h1;
  assign rom__T_755_data = 8'h0;
  assign rom__T_755_addr = 8'he6;
  assign rom__T_755_mask = 1'h1;
  assign rom__T_755_en = 1'h1;
  assign rom__T_758_data = 8'h0;
  assign rom__T_758_addr = 8'he7;
  assign rom__T_758_mask = 1'h1;
  assign rom__T_758_en = 1'h1;
  assign rom__T_762_data = 8'h0;
  assign rom__T_762_addr = 8'he8;
  assign rom__T_762_mask = 1'h1;
  assign rom__T_762_en = 1'h1;
  assign rom__T_765_data = 8'h0;
  assign rom__T_765_addr = 8'he9;
  assign rom__T_765_mask = 1'h1;
  assign rom__T_765_en = 1'h1;
  assign rom__T_768_data = 8'h0;
  assign rom__T_768_addr = 8'hea;
  assign rom__T_768_mask = 1'h1;
  assign rom__T_768_en = 1'h1;
  assign rom__T_771_data = 8'h0;
  assign rom__T_771_addr = 8'heb;
  assign rom__T_771_mask = 1'h1;
  assign rom__T_771_en = 1'h1;
  assign rom__T_775_data = 8'h0;
  assign rom__T_775_addr = 8'hec;
  assign rom__T_775_mask = 1'h1;
  assign rom__T_775_en = 1'h1;
  assign rom__T_778_data = 8'h0;
  assign rom__T_778_addr = 8'hed;
  assign rom__T_778_mask = 1'h1;
  assign rom__T_778_en = 1'h1;
  assign rom__T_781_data = 8'h0;
  assign rom__T_781_addr = 8'hee;
  assign rom__T_781_mask = 1'h1;
  assign rom__T_781_en = 1'h1;
  assign rom__T_784_data = 8'h0;
  assign rom__T_784_addr = 8'hef;
  assign rom__T_784_mask = 1'h1;
  assign rom__T_784_en = 1'h1;
  assign _T_787 = io_pc + 32'h3;
  assign _T_788 = _T_787[31:0];
  assign _T_789 = _T_788[7:0];
  assign _T_792 = io_pc + 32'h2;
  assign _T_793 = _T_792[31:0];
  assign _T_794 = _T_793[7:0];
  assign _T_797 = io_pc + 32'h1;
  assign _T_798 = _T_797[31:0];
  assign _T_799 = _T_798[7:0];
  assign _T_801 = io_pc[7:0];
  assign _T_803 = {rom__T_800_data,rom__T_802_data};
  assign _T_804 = {rom__T_790_data,rom__T_795_data};
  assign _T_805 = {_T_804,_T_803};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 240; initvar = initvar+1)
    rom[initvar] = _GEN_0[7:0];
  `endif
  _GEN_1 = {1{$random}};
  _GEN_2 = {1{$random}};
  _GEN_3 = {1{$random}};
  _GEN_4 = {1{$random}};
  end
`endif
  always @(posedge clock) begin
    if(rom__T_8_en & rom__T_8_mask) begin
      rom[rom__T_8_addr] <= rom__T_8_data;
    end
    if(rom__T_11_en & rom__T_11_mask) begin
      rom[rom__T_11_addr] <= rom__T_11_data;
    end
    if(rom__T_14_en & rom__T_14_mask) begin
      rom[rom__T_14_addr] <= rom__T_14_data;
    end
    if(rom__T_17_en & rom__T_17_mask) begin
      rom[rom__T_17_addr] <= rom__T_17_data;
    end
    if(rom__T_21_en & rom__T_21_mask) begin
      rom[rom__T_21_addr] <= rom__T_21_data;
    end
    if(rom__T_24_en & rom__T_24_mask) begin
      rom[rom__T_24_addr] <= rom__T_24_data;
    end
    if(rom__T_27_en & rom__T_27_mask) begin
      rom[rom__T_27_addr] <= rom__T_27_data;
    end
    if(rom__T_30_en & rom__T_30_mask) begin
      rom[rom__T_30_addr] <= rom__T_30_data;
    end
    if(rom__T_34_en & rom__T_34_mask) begin
      rom[rom__T_34_addr] <= rom__T_34_data;
    end
    if(rom__T_37_en & rom__T_37_mask) begin
      rom[rom__T_37_addr] <= rom__T_37_data;
    end
    if(rom__T_40_en & rom__T_40_mask) begin
      rom[rom__T_40_addr] <= rom__T_40_data;
    end
    if(rom__T_43_en & rom__T_43_mask) begin
      rom[rom__T_43_addr] <= rom__T_43_data;
    end
    if(rom__T_47_en & rom__T_47_mask) begin
      rom[rom__T_47_addr] <= rom__T_47_data;
    end
    if(rom__T_50_en & rom__T_50_mask) begin
      rom[rom__T_50_addr] <= rom__T_50_data;
    end
    if(rom__T_53_en & rom__T_53_mask) begin
      rom[rom__T_53_addr] <= rom__T_53_data;
    end
    if(rom__T_56_en & rom__T_56_mask) begin
      rom[rom__T_56_addr] <= rom__T_56_data;
    end
    if(rom__T_60_en & rom__T_60_mask) begin
      rom[rom__T_60_addr] <= rom__T_60_data;
    end
    if(rom__T_63_en & rom__T_63_mask) begin
      rom[rom__T_63_addr] <= rom__T_63_data;
    end
    if(rom__T_66_en & rom__T_66_mask) begin
      rom[rom__T_66_addr] <= rom__T_66_data;
    end
    if(rom__T_69_en & rom__T_69_mask) begin
      rom[rom__T_69_addr] <= rom__T_69_data;
    end
    if(rom__T_73_en & rom__T_73_mask) begin
      rom[rom__T_73_addr] <= rom__T_73_data;
    end
    if(rom__T_76_en & rom__T_76_mask) begin
      rom[rom__T_76_addr] <= rom__T_76_data;
    end
    if(rom__T_79_en & rom__T_79_mask) begin
      rom[rom__T_79_addr] <= rom__T_79_data;
    end
    if(rom__T_82_en & rom__T_82_mask) begin
      rom[rom__T_82_addr] <= rom__T_82_data;
    end
    if(rom__T_86_en & rom__T_86_mask) begin
      rom[rom__T_86_addr] <= rom__T_86_data;
    end
    if(rom__T_89_en & rom__T_89_mask) begin
      rom[rom__T_89_addr] <= rom__T_89_data;
    end
    if(rom__T_92_en & rom__T_92_mask) begin
      rom[rom__T_92_addr] <= rom__T_92_data;
    end
    if(rom__T_95_en & rom__T_95_mask) begin
      rom[rom__T_95_addr] <= rom__T_95_data;
    end
    if(rom__T_99_en & rom__T_99_mask) begin
      rom[rom__T_99_addr] <= rom__T_99_data;
    end
    if(rom__T_102_en & rom__T_102_mask) begin
      rom[rom__T_102_addr] <= rom__T_102_data;
    end
    if(rom__T_105_en & rom__T_105_mask) begin
      rom[rom__T_105_addr] <= rom__T_105_data;
    end
    if(rom__T_108_en & rom__T_108_mask) begin
      rom[rom__T_108_addr] <= rom__T_108_data;
    end
    if(rom__T_112_en & rom__T_112_mask) begin
      rom[rom__T_112_addr] <= rom__T_112_data;
    end
    if(rom__T_115_en & rom__T_115_mask) begin
      rom[rom__T_115_addr] <= rom__T_115_data;
    end
    if(rom__T_118_en & rom__T_118_mask) begin
      rom[rom__T_118_addr] <= rom__T_118_data;
    end
    if(rom__T_121_en & rom__T_121_mask) begin
      rom[rom__T_121_addr] <= rom__T_121_data;
    end
    if(rom__T_125_en & rom__T_125_mask) begin
      rom[rom__T_125_addr] <= rom__T_125_data;
    end
    if(rom__T_128_en & rom__T_128_mask) begin
      rom[rom__T_128_addr] <= rom__T_128_data;
    end
    if(rom__T_131_en & rom__T_131_mask) begin
      rom[rom__T_131_addr] <= rom__T_131_data;
    end
    if(rom__T_134_en & rom__T_134_mask) begin
      rom[rom__T_134_addr] <= rom__T_134_data;
    end
    if(rom__T_138_en & rom__T_138_mask) begin
      rom[rom__T_138_addr] <= rom__T_138_data;
    end
    if(rom__T_141_en & rom__T_141_mask) begin
      rom[rom__T_141_addr] <= rom__T_141_data;
    end
    if(rom__T_144_en & rom__T_144_mask) begin
      rom[rom__T_144_addr] <= rom__T_144_data;
    end
    if(rom__T_147_en & rom__T_147_mask) begin
      rom[rom__T_147_addr] <= rom__T_147_data;
    end
    if(rom__T_151_en & rom__T_151_mask) begin
      rom[rom__T_151_addr] <= rom__T_151_data;
    end
    if(rom__T_154_en & rom__T_154_mask) begin
      rom[rom__T_154_addr] <= rom__T_154_data;
    end
    if(rom__T_157_en & rom__T_157_mask) begin
      rom[rom__T_157_addr] <= rom__T_157_data;
    end
    if(rom__T_160_en & rom__T_160_mask) begin
      rom[rom__T_160_addr] <= rom__T_160_data;
    end
    if(rom__T_164_en & rom__T_164_mask) begin
      rom[rom__T_164_addr] <= rom__T_164_data;
    end
    if(rom__T_167_en & rom__T_167_mask) begin
      rom[rom__T_167_addr] <= rom__T_167_data;
    end
    if(rom__T_170_en & rom__T_170_mask) begin
      rom[rom__T_170_addr] <= rom__T_170_data;
    end
    if(rom__T_173_en & rom__T_173_mask) begin
      rom[rom__T_173_addr] <= rom__T_173_data;
    end
    if(rom__T_177_en & rom__T_177_mask) begin
      rom[rom__T_177_addr] <= rom__T_177_data;
    end
    if(rom__T_180_en & rom__T_180_mask) begin
      rom[rom__T_180_addr] <= rom__T_180_data;
    end
    if(rom__T_183_en & rom__T_183_mask) begin
      rom[rom__T_183_addr] <= rom__T_183_data;
    end
    if(rom__T_186_en & rom__T_186_mask) begin
      rom[rom__T_186_addr] <= rom__T_186_data;
    end
    if(rom__T_190_en & rom__T_190_mask) begin
      rom[rom__T_190_addr] <= rom__T_190_data;
    end
    if(rom__T_193_en & rom__T_193_mask) begin
      rom[rom__T_193_addr] <= rom__T_193_data;
    end
    if(rom__T_196_en & rom__T_196_mask) begin
      rom[rom__T_196_addr] <= rom__T_196_data;
    end
    if(rom__T_199_en & rom__T_199_mask) begin
      rom[rom__T_199_addr] <= rom__T_199_data;
    end
    if(rom__T_203_en & rom__T_203_mask) begin
      rom[rom__T_203_addr] <= rom__T_203_data;
    end
    if(rom__T_206_en & rom__T_206_mask) begin
      rom[rom__T_206_addr] <= rom__T_206_data;
    end
    if(rom__T_209_en & rom__T_209_mask) begin
      rom[rom__T_209_addr] <= rom__T_209_data;
    end
    if(rom__T_212_en & rom__T_212_mask) begin
      rom[rom__T_212_addr] <= rom__T_212_data;
    end
    if(rom__T_216_en & rom__T_216_mask) begin
      rom[rom__T_216_addr] <= rom__T_216_data;
    end
    if(rom__T_219_en & rom__T_219_mask) begin
      rom[rom__T_219_addr] <= rom__T_219_data;
    end
    if(rom__T_222_en & rom__T_222_mask) begin
      rom[rom__T_222_addr] <= rom__T_222_data;
    end
    if(rom__T_225_en & rom__T_225_mask) begin
      rom[rom__T_225_addr] <= rom__T_225_data;
    end
    if(rom__T_229_en & rom__T_229_mask) begin
      rom[rom__T_229_addr] <= rom__T_229_data;
    end
    if(rom__T_232_en & rom__T_232_mask) begin
      rom[rom__T_232_addr] <= rom__T_232_data;
    end
    if(rom__T_235_en & rom__T_235_mask) begin
      rom[rom__T_235_addr] <= rom__T_235_data;
    end
    if(rom__T_238_en & rom__T_238_mask) begin
      rom[rom__T_238_addr] <= rom__T_238_data;
    end
    if(rom__T_242_en & rom__T_242_mask) begin
      rom[rom__T_242_addr] <= rom__T_242_data;
    end
    if(rom__T_245_en & rom__T_245_mask) begin
      rom[rom__T_245_addr] <= rom__T_245_data;
    end
    if(rom__T_248_en & rom__T_248_mask) begin
      rom[rom__T_248_addr] <= rom__T_248_data;
    end
    if(rom__T_251_en & rom__T_251_mask) begin
      rom[rom__T_251_addr] <= rom__T_251_data;
    end
    if(rom__T_255_en & rom__T_255_mask) begin
      rom[rom__T_255_addr] <= rom__T_255_data;
    end
    if(rom__T_258_en & rom__T_258_mask) begin
      rom[rom__T_258_addr] <= rom__T_258_data;
    end
    if(rom__T_261_en & rom__T_261_mask) begin
      rom[rom__T_261_addr] <= rom__T_261_data;
    end
    if(rom__T_264_en & rom__T_264_mask) begin
      rom[rom__T_264_addr] <= rom__T_264_data;
    end
    if(rom__T_268_en & rom__T_268_mask) begin
      rom[rom__T_268_addr] <= rom__T_268_data;
    end
    if(rom__T_271_en & rom__T_271_mask) begin
      rom[rom__T_271_addr] <= rom__T_271_data;
    end
    if(rom__T_274_en & rom__T_274_mask) begin
      rom[rom__T_274_addr] <= rom__T_274_data;
    end
    if(rom__T_277_en & rom__T_277_mask) begin
      rom[rom__T_277_addr] <= rom__T_277_data;
    end
    if(rom__T_281_en & rom__T_281_mask) begin
      rom[rom__T_281_addr] <= rom__T_281_data;
    end
    if(rom__T_284_en & rom__T_284_mask) begin
      rom[rom__T_284_addr] <= rom__T_284_data;
    end
    if(rom__T_287_en & rom__T_287_mask) begin
      rom[rom__T_287_addr] <= rom__T_287_data;
    end
    if(rom__T_290_en & rom__T_290_mask) begin
      rom[rom__T_290_addr] <= rom__T_290_data;
    end
    if(rom__T_294_en & rom__T_294_mask) begin
      rom[rom__T_294_addr] <= rom__T_294_data;
    end
    if(rom__T_297_en & rom__T_297_mask) begin
      rom[rom__T_297_addr] <= rom__T_297_data;
    end
    if(rom__T_300_en & rom__T_300_mask) begin
      rom[rom__T_300_addr] <= rom__T_300_data;
    end
    if(rom__T_303_en & rom__T_303_mask) begin
      rom[rom__T_303_addr] <= rom__T_303_data;
    end
    if(rom__T_307_en & rom__T_307_mask) begin
      rom[rom__T_307_addr] <= rom__T_307_data;
    end
    if(rom__T_310_en & rom__T_310_mask) begin
      rom[rom__T_310_addr] <= rom__T_310_data;
    end
    if(rom__T_313_en & rom__T_313_mask) begin
      rom[rom__T_313_addr] <= rom__T_313_data;
    end
    if(rom__T_316_en & rom__T_316_mask) begin
      rom[rom__T_316_addr] <= rom__T_316_data;
    end
    if(rom__T_320_en & rom__T_320_mask) begin
      rom[rom__T_320_addr] <= rom__T_320_data;
    end
    if(rom__T_323_en & rom__T_323_mask) begin
      rom[rom__T_323_addr] <= rom__T_323_data;
    end
    if(rom__T_326_en & rom__T_326_mask) begin
      rom[rom__T_326_addr] <= rom__T_326_data;
    end
    if(rom__T_329_en & rom__T_329_mask) begin
      rom[rom__T_329_addr] <= rom__T_329_data;
    end
    if(rom__T_333_en & rom__T_333_mask) begin
      rom[rom__T_333_addr] <= rom__T_333_data;
    end
    if(rom__T_336_en & rom__T_336_mask) begin
      rom[rom__T_336_addr] <= rom__T_336_data;
    end
    if(rom__T_339_en & rom__T_339_mask) begin
      rom[rom__T_339_addr] <= rom__T_339_data;
    end
    if(rom__T_342_en & rom__T_342_mask) begin
      rom[rom__T_342_addr] <= rom__T_342_data;
    end
    if(rom__T_346_en & rom__T_346_mask) begin
      rom[rom__T_346_addr] <= rom__T_346_data;
    end
    if(rom__T_349_en & rom__T_349_mask) begin
      rom[rom__T_349_addr] <= rom__T_349_data;
    end
    if(rom__T_352_en & rom__T_352_mask) begin
      rom[rom__T_352_addr] <= rom__T_352_data;
    end
    if(rom__T_355_en & rom__T_355_mask) begin
      rom[rom__T_355_addr] <= rom__T_355_data;
    end
    if(rom__T_359_en & rom__T_359_mask) begin
      rom[rom__T_359_addr] <= rom__T_359_data;
    end
    if(rom__T_362_en & rom__T_362_mask) begin
      rom[rom__T_362_addr] <= rom__T_362_data;
    end
    if(rom__T_365_en & rom__T_365_mask) begin
      rom[rom__T_365_addr] <= rom__T_365_data;
    end
    if(rom__T_368_en & rom__T_368_mask) begin
      rom[rom__T_368_addr] <= rom__T_368_data;
    end
    if(rom__T_372_en & rom__T_372_mask) begin
      rom[rom__T_372_addr] <= rom__T_372_data;
    end
    if(rom__T_375_en & rom__T_375_mask) begin
      rom[rom__T_375_addr] <= rom__T_375_data;
    end
    if(rom__T_378_en & rom__T_378_mask) begin
      rom[rom__T_378_addr] <= rom__T_378_data;
    end
    if(rom__T_381_en & rom__T_381_mask) begin
      rom[rom__T_381_addr] <= rom__T_381_data;
    end
    if(rom__T_385_en & rom__T_385_mask) begin
      rom[rom__T_385_addr] <= rom__T_385_data;
    end
    if(rom__T_388_en & rom__T_388_mask) begin
      rom[rom__T_388_addr] <= rom__T_388_data;
    end
    if(rom__T_391_en & rom__T_391_mask) begin
      rom[rom__T_391_addr] <= rom__T_391_data;
    end
    if(rom__T_394_en & rom__T_394_mask) begin
      rom[rom__T_394_addr] <= rom__T_394_data;
    end
    if(rom__T_398_en & rom__T_398_mask) begin
      rom[rom__T_398_addr] <= rom__T_398_data;
    end
    if(rom__T_401_en & rom__T_401_mask) begin
      rom[rom__T_401_addr] <= rom__T_401_data;
    end
    if(rom__T_404_en & rom__T_404_mask) begin
      rom[rom__T_404_addr] <= rom__T_404_data;
    end
    if(rom__T_407_en & rom__T_407_mask) begin
      rom[rom__T_407_addr] <= rom__T_407_data;
    end
    if(rom__T_411_en & rom__T_411_mask) begin
      rom[rom__T_411_addr] <= rom__T_411_data;
    end
    if(rom__T_414_en & rom__T_414_mask) begin
      rom[rom__T_414_addr] <= rom__T_414_data;
    end
    if(rom__T_417_en & rom__T_417_mask) begin
      rom[rom__T_417_addr] <= rom__T_417_data;
    end
    if(rom__T_420_en & rom__T_420_mask) begin
      rom[rom__T_420_addr] <= rom__T_420_data;
    end
    if(rom__T_424_en & rom__T_424_mask) begin
      rom[rom__T_424_addr] <= rom__T_424_data;
    end
    if(rom__T_427_en & rom__T_427_mask) begin
      rom[rom__T_427_addr] <= rom__T_427_data;
    end
    if(rom__T_430_en & rom__T_430_mask) begin
      rom[rom__T_430_addr] <= rom__T_430_data;
    end
    if(rom__T_433_en & rom__T_433_mask) begin
      rom[rom__T_433_addr] <= rom__T_433_data;
    end
    if(rom__T_437_en & rom__T_437_mask) begin
      rom[rom__T_437_addr] <= rom__T_437_data;
    end
    if(rom__T_440_en & rom__T_440_mask) begin
      rom[rom__T_440_addr] <= rom__T_440_data;
    end
    if(rom__T_443_en & rom__T_443_mask) begin
      rom[rom__T_443_addr] <= rom__T_443_data;
    end
    if(rom__T_446_en & rom__T_446_mask) begin
      rom[rom__T_446_addr] <= rom__T_446_data;
    end
    if(rom__T_450_en & rom__T_450_mask) begin
      rom[rom__T_450_addr] <= rom__T_450_data;
    end
    if(rom__T_453_en & rom__T_453_mask) begin
      rom[rom__T_453_addr] <= rom__T_453_data;
    end
    if(rom__T_456_en & rom__T_456_mask) begin
      rom[rom__T_456_addr] <= rom__T_456_data;
    end
    if(rom__T_459_en & rom__T_459_mask) begin
      rom[rom__T_459_addr] <= rom__T_459_data;
    end
    if(rom__T_463_en & rom__T_463_mask) begin
      rom[rom__T_463_addr] <= rom__T_463_data;
    end
    if(rom__T_466_en & rom__T_466_mask) begin
      rom[rom__T_466_addr] <= rom__T_466_data;
    end
    if(rom__T_469_en & rom__T_469_mask) begin
      rom[rom__T_469_addr] <= rom__T_469_data;
    end
    if(rom__T_472_en & rom__T_472_mask) begin
      rom[rom__T_472_addr] <= rom__T_472_data;
    end
    if(rom__T_476_en & rom__T_476_mask) begin
      rom[rom__T_476_addr] <= rom__T_476_data;
    end
    if(rom__T_479_en & rom__T_479_mask) begin
      rom[rom__T_479_addr] <= rom__T_479_data;
    end
    if(rom__T_482_en & rom__T_482_mask) begin
      rom[rom__T_482_addr] <= rom__T_482_data;
    end
    if(rom__T_485_en & rom__T_485_mask) begin
      rom[rom__T_485_addr] <= rom__T_485_data;
    end
    if(rom__T_489_en & rom__T_489_mask) begin
      rom[rom__T_489_addr] <= rom__T_489_data;
    end
    if(rom__T_492_en & rom__T_492_mask) begin
      rom[rom__T_492_addr] <= rom__T_492_data;
    end
    if(rom__T_495_en & rom__T_495_mask) begin
      rom[rom__T_495_addr] <= rom__T_495_data;
    end
    if(rom__T_498_en & rom__T_498_mask) begin
      rom[rom__T_498_addr] <= rom__T_498_data;
    end
    if(rom__T_502_en & rom__T_502_mask) begin
      rom[rom__T_502_addr] <= rom__T_502_data;
    end
    if(rom__T_505_en & rom__T_505_mask) begin
      rom[rom__T_505_addr] <= rom__T_505_data;
    end
    if(rom__T_508_en & rom__T_508_mask) begin
      rom[rom__T_508_addr] <= rom__T_508_data;
    end
    if(rom__T_511_en & rom__T_511_mask) begin
      rom[rom__T_511_addr] <= rom__T_511_data;
    end
    if(rom__T_515_en & rom__T_515_mask) begin
      rom[rom__T_515_addr] <= rom__T_515_data;
    end
    if(rom__T_518_en & rom__T_518_mask) begin
      rom[rom__T_518_addr] <= rom__T_518_data;
    end
    if(rom__T_521_en & rom__T_521_mask) begin
      rom[rom__T_521_addr] <= rom__T_521_data;
    end
    if(rom__T_524_en & rom__T_524_mask) begin
      rom[rom__T_524_addr] <= rom__T_524_data;
    end
    if(rom__T_528_en & rom__T_528_mask) begin
      rom[rom__T_528_addr] <= rom__T_528_data;
    end
    if(rom__T_531_en & rom__T_531_mask) begin
      rom[rom__T_531_addr] <= rom__T_531_data;
    end
    if(rom__T_534_en & rom__T_534_mask) begin
      rom[rom__T_534_addr] <= rom__T_534_data;
    end
    if(rom__T_537_en & rom__T_537_mask) begin
      rom[rom__T_537_addr] <= rom__T_537_data;
    end
    if(rom__T_541_en & rom__T_541_mask) begin
      rom[rom__T_541_addr] <= rom__T_541_data;
    end
    if(rom__T_544_en & rom__T_544_mask) begin
      rom[rom__T_544_addr] <= rom__T_544_data;
    end
    if(rom__T_547_en & rom__T_547_mask) begin
      rom[rom__T_547_addr] <= rom__T_547_data;
    end
    if(rom__T_550_en & rom__T_550_mask) begin
      rom[rom__T_550_addr] <= rom__T_550_data;
    end
    if(rom__T_554_en & rom__T_554_mask) begin
      rom[rom__T_554_addr] <= rom__T_554_data;
    end
    if(rom__T_557_en & rom__T_557_mask) begin
      rom[rom__T_557_addr] <= rom__T_557_data;
    end
    if(rom__T_560_en & rom__T_560_mask) begin
      rom[rom__T_560_addr] <= rom__T_560_data;
    end
    if(rom__T_563_en & rom__T_563_mask) begin
      rom[rom__T_563_addr] <= rom__T_563_data;
    end
    if(rom__T_567_en & rom__T_567_mask) begin
      rom[rom__T_567_addr] <= rom__T_567_data;
    end
    if(rom__T_570_en & rom__T_570_mask) begin
      rom[rom__T_570_addr] <= rom__T_570_data;
    end
    if(rom__T_573_en & rom__T_573_mask) begin
      rom[rom__T_573_addr] <= rom__T_573_data;
    end
    if(rom__T_576_en & rom__T_576_mask) begin
      rom[rom__T_576_addr] <= rom__T_576_data;
    end
    if(rom__T_580_en & rom__T_580_mask) begin
      rom[rom__T_580_addr] <= rom__T_580_data;
    end
    if(rom__T_583_en & rom__T_583_mask) begin
      rom[rom__T_583_addr] <= rom__T_583_data;
    end
    if(rom__T_586_en & rom__T_586_mask) begin
      rom[rom__T_586_addr] <= rom__T_586_data;
    end
    if(rom__T_589_en & rom__T_589_mask) begin
      rom[rom__T_589_addr] <= rom__T_589_data;
    end
    if(rom__T_593_en & rom__T_593_mask) begin
      rom[rom__T_593_addr] <= rom__T_593_data;
    end
    if(rom__T_596_en & rom__T_596_mask) begin
      rom[rom__T_596_addr] <= rom__T_596_data;
    end
    if(rom__T_599_en & rom__T_599_mask) begin
      rom[rom__T_599_addr] <= rom__T_599_data;
    end
    if(rom__T_602_en & rom__T_602_mask) begin
      rom[rom__T_602_addr] <= rom__T_602_data;
    end
    if(rom__T_606_en & rom__T_606_mask) begin
      rom[rom__T_606_addr] <= rom__T_606_data;
    end
    if(rom__T_609_en & rom__T_609_mask) begin
      rom[rom__T_609_addr] <= rom__T_609_data;
    end
    if(rom__T_612_en & rom__T_612_mask) begin
      rom[rom__T_612_addr] <= rom__T_612_data;
    end
    if(rom__T_615_en & rom__T_615_mask) begin
      rom[rom__T_615_addr] <= rom__T_615_data;
    end
    if(rom__T_619_en & rom__T_619_mask) begin
      rom[rom__T_619_addr] <= rom__T_619_data;
    end
    if(rom__T_622_en & rom__T_622_mask) begin
      rom[rom__T_622_addr] <= rom__T_622_data;
    end
    if(rom__T_625_en & rom__T_625_mask) begin
      rom[rom__T_625_addr] <= rom__T_625_data;
    end
    if(rom__T_628_en & rom__T_628_mask) begin
      rom[rom__T_628_addr] <= rom__T_628_data;
    end
    if(rom__T_632_en & rom__T_632_mask) begin
      rom[rom__T_632_addr] <= rom__T_632_data;
    end
    if(rom__T_635_en & rom__T_635_mask) begin
      rom[rom__T_635_addr] <= rom__T_635_data;
    end
    if(rom__T_638_en & rom__T_638_mask) begin
      rom[rom__T_638_addr] <= rom__T_638_data;
    end
    if(rom__T_641_en & rom__T_641_mask) begin
      rom[rom__T_641_addr] <= rom__T_641_data;
    end
    if(rom__T_645_en & rom__T_645_mask) begin
      rom[rom__T_645_addr] <= rom__T_645_data;
    end
    if(rom__T_648_en & rom__T_648_mask) begin
      rom[rom__T_648_addr] <= rom__T_648_data;
    end
    if(rom__T_651_en & rom__T_651_mask) begin
      rom[rom__T_651_addr] <= rom__T_651_data;
    end
    if(rom__T_654_en & rom__T_654_mask) begin
      rom[rom__T_654_addr] <= rom__T_654_data;
    end
    if(rom__T_658_en & rom__T_658_mask) begin
      rom[rom__T_658_addr] <= rom__T_658_data;
    end
    if(rom__T_661_en & rom__T_661_mask) begin
      rom[rom__T_661_addr] <= rom__T_661_data;
    end
    if(rom__T_664_en & rom__T_664_mask) begin
      rom[rom__T_664_addr] <= rom__T_664_data;
    end
    if(rom__T_667_en & rom__T_667_mask) begin
      rom[rom__T_667_addr] <= rom__T_667_data;
    end
    if(rom__T_671_en & rom__T_671_mask) begin
      rom[rom__T_671_addr] <= rom__T_671_data;
    end
    if(rom__T_674_en & rom__T_674_mask) begin
      rom[rom__T_674_addr] <= rom__T_674_data;
    end
    if(rom__T_677_en & rom__T_677_mask) begin
      rom[rom__T_677_addr] <= rom__T_677_data;
    end
    if(rom__T_680_en & rom__T_680_mask) begin
      rom[rom__T_680_addr] <= rom__T_680_data;
    end
    if(rom__T_684_en & rom__T_684_mask) begin
      rom[rom__T_684_addr] <= rom__T_684_data;
    end
    if(rom__T_687_en & rom__T_687_mask) begin
      rom[rom__T_687_addr] <= rom__T_687_data;
    end
    if(rom__T_690_en & rom__T_690_mask) begin
      rom[rom__T_690_addr] <= rom__T_690_data;
    end
    if(rom__T_693_en & rom__T_693_mask) begin
      rom[rom__T_693_addr] <= rom__T_693_data;
    end
    if(rom__T_697_en & rom__T_697_mask) begin
      rom[rom__T_697_addr] <= rom__T_697_data;
    end
    if(rom__T_700_en & rom__T_700_mask) begin
      rom[rom__T_700_addr] <= rom__T_700_data;
    end
    if(rom__T_703_en & rom__T_703_mask) begin
      rom[rom__T_703_addr] <= rom__T_703_data;
    end
    if(rom__T_706_en & rom__T_706_mask) begin
      rom[rom__T_706_addr] <= rom__T_706_data;
    end
    if(rom__T_710_en & rom__T_710_mask) begin
      rom[rom__T_710_addr] <= rom__T_710_data;
    end
    if(rom__T_713_en & rom__T_713_mask) begin
      rom[rom__T_713_addr] <= rom__T_713_data;
    end
    if(rom__T_716_en & rom__T_716_mask) begin
      rom[rom__T_716_addr] <= rom__T_716_data;
    end
    if(rom__T_719_en & rom__T_719_mask) begin
      rom[rom__T_719_addr] <= rom__T_719_data;
    end
    if(rom__T_723_en & rom__T_723_mask) begin
      rom[rom__T_723_addr] <= rom__T_723_data;
    end
    if(rom__T_726_en & rom__T_726_mask) begin
      rom[rom__T_726_addr] <= rom__T_726_data;
    end
    if(rom__T_729_en & rom__T_729_mask) begin
      rom[rom__T_729_addr] <= rom__T_729_data;
    end
    if(rom__T_732_en & rom__T_732_mask) begin
      rom[rom__T_732_addr] <= rom__T_732_data;
    end
    if(rom__T_736_en & rom__T_736_mask) begin
      rom[rom__T_736_addr] <= rom__T_736_data;
    end
    if(rom__T_739_en & rom__T_739_mask) begin
      rom[rom__T_739_addr] <= rom__T_739_data;
    end
    if(rom__T_742_en & rom__T_742_mask) begin
      rom[rom__T_742_addr] <= rom__T_742_data;
    end
    if(rom__T_745_en & rom__T_745_mask) begin
      rom[rom__T_745_addr] <= rom__T_745_data;
    end
    if(rom__T_749_en & rom__T_749_mask) begin
      rom[rom__T_749_addr] <= rom__T_749_data;
    end
    if(rom__T_752_en & rom__T_752_mask) begin
      rom[rom__T_752_addr] <= rom__T_752_data;
    end
    if(rom__T_755_en & rom__T_755_mask) begin
      rom[rom__T_755_addr] <= rom__T_755_data;
    end
    if(rom__T_758_en & rom__T_758_mask) begin
      rom[rom__T_758_addr] <= rom__T_758_data;
    end
    if(rom__T_762_en & rom__T_762_mask) begin
      rom[rom__T_762_addr] <= rom__T_762_data;
    end
    if(rom__T_765_en & rom__T_765_mask) begin
      rom[rom__T_765_addr] <= rom__T_765_data;
    end
    if(rom__T_768_en & rom__T_768_mask) begin
      rom[rom__T_768_addr] <= rom__T_768_data;
    end
    if(rom__T_771_en & rom__T_771_mask) begin
      rom[rom__T_771_addr] <= rom__T_771_data;
    end
    if(rom__T_775_en & rom__T_775_mask) begin
      rom[rom__T_775_addr] <= rom__T_775_data;
    end
    if(rom__T_778_en & rom__T_778_mask) begin
      rom[rom__T_778_addr] <= rom__T_778_data;
    end
    if(rom__T_781_en & rom__T_781_mask) begin
      rom[rom__T_781_addr] <= rom__T_781_data;
    end
    if(rom__T_784_en & rom__T_784_mask) begin
      rom[rom__T_784_addr] <= rom__T_784_data;
    end
  end
endmodule
module ProgramCounter(
  input         clock,
  input         reset,
  input         io_branch,
  input  [31:0] io_pc_src,
  output [31:0] io_pc_next,
  output [31:0] io_pc
);
  reg [31:0] pc_reg;
  reg [31:0] _GEN_0;
  wire [32:0] _T_8;
  wire [31:0] _T_9;
  wire [31:0] _T_10;
  assign io_pc_next = _T_9;
  assign io_pc = pc_reg;
  assign _T_8 = pc_reg + 32'h4;
  assign _T_9 = _T_8[31:0];
  assign _T_10 = io_branch ? io_pc_src : io_pc_next;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_0 = {1{$random}};
  pc_reg = _GEN_0[31:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (reset) begin
      pc_reg <= 32'h54;
    end else begin
      if (io_branch) begin
        pc_reg <= io_pc_src;
      end else begin
        pc_reg <= io_pc_next;
      end
    end
  end
endmodule
module Decoder(
  input  [31:0] io_inst,
  output [6:0]  io_ctrl_opcode,
  output [2:0]  io_ctrl_funct3,
  output [6:0]  io_ctrl_funct7,
  output [4:0]  io_rs_rs1,
  output [4:0]  io_rs_rs2,
  output [4:0]  io_rd,
  output [31:0] io_imm
);
  wire [6:0] _T_17;
  wire [4:0] _T_18;
  wire [2:0] _T_19;
  wire [4:0] _T_20;
  wire [4:0] _T_21;
  wire  _T_22;
  wire [6:0] _T_23;
  wire [6:0] _T_25;
  wire [11:0] _T_28;
  wire [31:0] _T_29;
  wire  _T_30;
  wire [31:0] _GEN_1;
  wire  _T_34;
  wire [31:0] _GEN_2;
  wire  _T_38;
  wire [26:0] _T_42;
  wire [31:0] _T_43;
  wire [31:0] _GEN_3;
  wire  _T_44;
  wire  _T_46;
  wire  _T_47;
  wire [5:0] _T_48;
  wire [3:0] _T_49;
  wire [9:0] _T_50;
  wire [20:0] _T_51;
  wire [21:0] _T_52;
  wire [31:0] _T_53;
  wire [31:0] _GEN_4;
  wire  _T_54;
  wire [19:0] _T_56;
  wire [31:0] _T_57;
  wire [31:0] _GEN_5;
  wire  _T_58;
  wire [31:0] _GEN_6;
  wire  _T_62;
  wire [7:0] _T_65;
  wire  _T_66;
  wire [9:0] _T_67;
  wire [10:0] _T_69;
  wire [11:0] _T_70;
  wire [11:0] _T_71;
  wire [19:0] _T_72;
  wire [31:0] _T_73;
  wire [31:0] _GEN_7;
  assign io_ctrl_opcode = _T_17;
  assign io_ctrl_funct3 = _T_19;
  assign io_ctrl_funct7 = _T_25;
  assign io_rs_rs1 = _T_20;
  assign io_rs_rs2 = _T_21;
  assign io_rd = _T_18;
  assign io_imm = _GEN_7;
  assign _T_17 = io_inst[6:0];
  assign _T_18 = io_inst[11:7];
  assign _T_19 = io_inst[14:12];
  assign _T_20 = io_inst[19:15];
  assign _T_21 = io_inst[24:20];
  assign _T_22 = io_ctrl_opcode == 7'h33;
  assign _T_23 = io_inst[31:25];
  assign _T_25 = _T_22 ? _T_23 : 7'h0;
  assign _T_28 = io_inst[31:20];
  assign _T_29 = {20'h0,_T_28};
  assign _T_30 = 7'h3 == io_ctrl_opcode;
  assign _GEN_1 = _T_30 ? _T_29 : _T_29;
  assign _T_34 = 7'h67 == io_ctrl_opcode;
  assign _GEN_2 = _T_34 ? _T_29 : _GEN_1;
  assign _T_38 = 7'h23 == io_ctrl_opcode;
  assign _T_42 = {20'h0,_T_23};
  assign _T_43 = {_T_42,_T_18};
  assign _GEN_3 = _T_38 ? _T_43 : _GEN_2;
  assign _T_44 = 7'h63 == io_ctrl_opcode;
  assign _T_46 = io_inst[31];
  assign _T_47 = io_inst[7];
  assign _T_48 = io_inst[30:25];
  assign _T_49 = io_inst[11:8];
  assign _T_50 = {_T_48,_T_49};
  assign _T_51 = {20'h0,_T_46};
  assign _T_52 = {_T_51,_T_47};
  assign _T_53 = {_T_52,_T_50};
  assign _GEN_4 = _T_44 ? _T_53 : _GEN_3;
  assign _T_54 = 7'h37 == io_ctrl_opcode;
  assign _T_56 = io_inst[31:12];
  assign _T_57 = {12'h0,_T_56};
  assign _GEN_5 = _T_54 ? _T_57 : _GEN_4;
  assign _T_58 = 7'h17 == io_ctrl_opcode;
  assign _GEN_6 = _T_58 ? _T_57 : _GEN_5;
  assign _T_62 = 7'h6f == io_ctrl_opcode;
  assign _T_65 = io_inst[19:12];
  assign _T_66 = io_inst[20];
  assign _T_67 = io_inst[30:21];
  assign _T_69 = {_T_66,_T_67};
  assign _T_70 = {_T_69,1'h0};
  assign _T_71 = {11'h0,_T_46};
  assign _T_72 = {_T_71,_T_65};
  assign _T_73 = {_T_72,_T_70};
  assign _GEN_7 = _T_62 ? _T_73 : _GEN_6;
endmodule
module Control(
  input  [6:0] io_ctrl_opcode,
  input  [2:0] io_ctrl_funct3,
  input  [6:0] io_ctrl_funct7,
  output       io_WB_reg_w,
  output       io_WB_rd_mem,
  output       io_MEM_branch,
  output       io_MEM_write,
  output       io_MEM_read,
  output [2:0] io_MEM_func,
  output [6:0] io_EX_opcode,
  output       io_EX_alu_sel,
  output       io_EX_dst_sel,
  output [2:0] io_EX_alu_op_func,
  output       io_EX_alu_op_alt
);
  wire  _T_30;
  wire  _T_31;
  wire  _T_32;
  wire  _T_33;
  wire  _T_34;
  wire  _T_35;
  wire  _T_36;
  wire  _T_37;
  wire  _T_38;
  wire  _T_39;
  wire  _T_41;
  assign io_WB_reg_w = _T_41;
  assign io_WB_rd_mem = io_MEM_read;
  assign io_MEM_branch = _T_36;
  assign io_MEM_write = _T_35;
  assign io_MEM_read = _T_34;
  assign io_MEM_func = io_ctrl_funct3;
  assign io_EX_opcode = io_ctrl_opcode;
  assign io_EX_alu_sel = _T_30;
  assign io_EX_dst_sel = _T_31;
  assign io_EX_alu_op_func = io_ctrl_funct3;
  assign io_EX_alu_op_alt = _T_33;
  assign _T_30 = io_ctrl_opcode != 7'h33;
  assign _T_31 = io_ctrl_opcode != 7'h3;
  assign _T_32 = io_ctrl_funct7[5];
  assign _T_33 = io_EX_alu_sel ? 1'h0 : _T_32;
  assign _T_34 = io_ctrl_opcode == 7'h3;
  assign _T_35 = io_ctrl_opcode == 7'h23;
  assign _T_36 = io_ctrl_opcode == 7'h63;
  assign _T_37 = io_ctrl_opcode == 7'h33;
  assign _T_38 = io_ctrl_opcode == 7'h13;
  assign _T_39 = _T_37 | _T_38;
  assign _T_41 = _T_39 | _T_34;
endmodule
module Registers(
  input         clock,
  input  [4:0]  io_rs_rs1,
  input  [4:0]  io_rs_rs2,
  input         io_reg_w,
  input  [4:0]  io_rd,
  input  [31:0] io_res,
  output [31:0] io_op_op1,
  output [31:0] io_op_op2
);
  reg [31:0] x [0:31];
  reg [31:0] _GEN_0;
  wire [31:0] x__T_23_data;
  wire [4:0] x__T_23_addr;
  wire [31:0] x__T_25_data;
  wire [4:0] x__T_25_addr;
  wire [31:0] x__T_15_data;
  wire [4:0] x__T_15_addr;
  wire  x__T_15_mask;
  wire  x__T_15_en;
  wire [31:0] x__T_16_data;
  wire [4:0] x__T_16_addr;
  wire  x__T_16_mask;
  wire  x__T_16_en;
  wire  _T_17;
  wire  _T_18;
  wire  _T_19;
  wire  fwd_rs1;
  wire  _T_22;
  wire  fwd_rs2;
  wire [31:0] _T_24;
  wire [31:0] _T_26;
  assign io_op_op1 = _T_24;
  assign io_op_op2 = _T_26;
  assign x__T_23_addr = io_rs_rs1;
  assign x__T_23_data = x[x__T_23_addr];
  assign x__T_25_addr = io_rs_rs2;
  assign x__T_25_data = x[x__T_25_addr];
  assign x__T_15_data = 32'h0;
  assign x__T_15_addr = 5'h0;
  assign x__T_15_mask = 1'h1;
  assign x__T_15_en = 1'h1;
  assign x__T_16_data = io_res;
  assign x__T_16_addr = io_rd;
  assign x__T_16_mask = io_reg_w;
  assign x__T_16_en = io_reg_w;
  assign _T_17 = io_res != 32'h0;
  assign _T_18 = io_reg_w & _T_17;
  assign _T_19 = io_rd == io_rs_rs1;
  assign fwd_rs1 = _T_18 & _T_19;
  assign _T_22 = io_rd == io_rs_rs2;
  assign fwd_rs2 = _T_18 & _T_22;
  assign _T_24 = fwd_rs1 ? io_res : x__T_23_data;
  assign _T_26 = fwd_rs2 ? io_res : x__T_25_data;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    x[initvar] = _GEN_0[31:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if(x__T_15_en & x__T_15_mask) begin
      x[x__T_15_addr] <= x__T_15_data;
    end
    if(x__T_16_en & x__T_16_mask) begin
      x[x__T_16_addr] <= x__T_16_data;
    end
  end
endmodule
module ALU(
  input  [6:0]  io_opcode,
  input  [2:0]  io_alu_op_func,
  input         io_alu_op_alt,
  input  [31:0] io_op_op1,
  input  [31:0] io_op_op2,
  output [31:0] io_res
);
  wire [4:0] shamt;
  wire [32:0] _T_10;
  wire [32:0] _T_11;
  wire [31:0] _T_12;
  wire [32:0] _T_13;
  wire [31:0] _T_14;
  wire [31:0] _T_15;
  wire [62:0] _GEN_0;
  wire [62:0] _T_16;
  wire  _T_17;
  wire [31:0] _T_18;
  wire [31:0] _T_19;
  wire [31:0] _T_20;
  wire [31:0] _T_21;
  wire  _T_22;
  wire [31:0] _T_23;
  wire  _T_24;
  wire [31:0] _T_25;
  wire  _T_26;
  wire [31:0] _T_27;
  wire  _T_28;
  wire [31:0] _T_29;
  wire  _T_30;
  wire [62:0] _T_31;
  wire  _T_32;
  wire [62:0] _T_33;
  wire [62:0] _T_53;
  wire  _T_61;
  wire [31:0] _T_62;
  wire  _T_63;
  wire [31:0] _T_64;
  wire  _T_65;
  wire [31:0] _T_66;
  wire  _T_67;
  wire [62:0] _T_68;
  wire  _T_69;
  wire [62:0] _T_70;
  reg  _GEN_1;
  reg [31:0] _GEN_2;
  assign io_res = _T_70[31:0];
  assign shamt = io_op_op2[4:0];
  assign _T_10 = io_op_op1 - io_op_op2;
  assign _T_11 = $unsigned(_T_10);
  assign _T_12 = _T_11[31:0];
  assign _T_13 = io_op_op1 + io_op_op2;
  assign _T_14 = _T_13[31:0];
  assign _T_15 = io_alu_op_alt ? _T_12 : _T_14;
  assign _GEN_0 = {{31'd0}, io_op_op1};
  assign _T_16 = _GEN_0 << shamt;
  assign _T_17 = io_op_op1 < io_op_op2;
  assign _T_18 = io_op_op1 ^ io_op_op2;
  assign _T_19 = io_op_op1 >> shamt;
  assign _T_20 = io_alu_op_alt ? 32'h0 : _T_19;
  assign _T_21 = io_op_op1 | io_op_op2;
  assign _T_22 = 3'h6 == io_alu_op_func;
  assign _T_23 = _T_22 ? _T_21 : 32'h0;
  assign _T_24 = 3'h5 == io_alu_op_func;
  assign _T_25 = _T_24 ? _T_20 : _T_23;
  assign _T_26 = 3'h4 == io_alu_op_func;
  assign _T_27 = _T_26 ? _T_18 : _T_25;
  assign _T_28 = 3'h3 == io_alu_op_func;
  assign _T_29 = _T_28 ? {{31'd0}, _T_17} : _T_27;
  assign _T_30 = 3'h1 == io_alu_op_func;
  assign _T_31 = _T_30 ? _T_16 : {{31'd0}, _T_29};
  assign _T_32 = 3'h0 == io_alu_op_func;
  assign _T_33 = _T_32 ? {{31'd0}, _T_15} : _T_31;
  assign _T_53 = _T_32 ? {{31'd0}, _T_14} : _T_31;
  assign _T_61 = 7'h63 == io_opcode;
  assign _T_62 = _T_61 ? _T_12 : 32'h0;
  assign _T_63 = 7'h23 == io_opcode;
  assign _T_64 = _T_63 ? _T_14 : _T_62;
  assign _T_65 = 7'h3 == io_opcode;
  assign _T_66 = _T_65 ? _T_14 : _T_64;
  assign _T_67 = 7'h13 == io_opcode;
  assign _T_68 = _T_67 ? _T_53 : {{31'd0}, _T_66};
  assign _T_69 = 7'h33 == io_opcode;
  assign _T_70 = _T_69 ? _T_33 : _T_68;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2 = {1{$random}};
  _GEN_1 = _GEN_2[0:0];
  `endif
  end
`endif
endmodule
module DataMemory(
  input         clock,
  input         io_mem_write,
  input         io_mem_read,
  input  [2:0]  io_mem_func,
  input  [31:0] io_op_op1,
  input  [31:0] io_op_op2,
  output [31:0] io_res
);
  reg [7:0] data_mem [0:511];
  reg [31:0] _GEN_0;
  wire [7:0] data_mem__T_49_data;
  wire [8:0] data_mem__T_49_addr;
  wire [7:0] data_mem__T_55_data;
  wire [8:0] data_mem__T_55_addr;
  wire [7:0] data_mem__T_57_data;
  wire [8:0] data_mem__T_57_addr;
  wire [7:0] data_mem__T_64_data;
  wire [8:0] data_mem__T_64_addr;
  wire [7:0] data_mem__T_69_data;
  wire [8:0] data_mem__T_69_addr;
  wire [7:0] data_mem__T_74_data;
  wire [8:0] data_mem__T_74_addr;
  wire [7:0] data_mem__T_76_data;
  wire [8:0] data_mem__T_76_addr;
  wire [7:0] data_mem__T_13_data;
  wire [8:0] data_mem__T_13_addr;
  wire  data_mem__T_13_mask;
  wire  data_mem__T_13_en;
  wire [7:0] data_mem__T_17_data;
  wire [8:0] data_mem__T_17_addr;
  wire  data_mem__T_17_mask;
  wire  data_mem__T_17_en;
  wire [7:0] data_mem__T_23_data;
  wire [8:0] data_mem__T_23_addr;
  wire  data_mem__T_23_mask;
  wire  data_mem__T_23_en;
  wire [7:0] data_mem__T_27_data;
  wire [8:0] data_mem__T_27_addr;
  wire  data_mem__T_27_mask;
  wire  data_mem__T_27_en;
  wire [7:0] data_mem__T_33_data;
  wire [8:0] data_mem__T_33_addr;
  wire  data_mem__T_33_mask;
  wire  data_mem__T_33_en;
  wire [7:0] data_mem__T_39_data;
  wire [8:0] data_mem__T_39_addr;
  wire  data_mem__T_39_mask;
  wire  data_mem__T_39_en;
  wire [7:0] data_mem__T_45_data;
  wire [8:0] data_mem__T_45_addr;
  wire  data_mem__T_45_mask;
  wire  data_mem__T_45_en;
  wire  _T_11;
  wire [8:0] _T_12;
  wire [7:0] _T_14;
  wire  _T_15;
  wire [8:0] _T_16;
  wire [7:0] _T_18;
  wire [32:0] _T_20;
  wire [31:0] _T_21;
  wire [8:0] _T_22;
  wire [7:0] _T_24;
  wire  _T_25;
  wire [8:0] _T_26;
  wire [7:0] _T_28;
  wire [8:0] _T_32;
  wire [7:0] _T_34;
  wire [32:0] _T_36;
  wire [31:0] _T_37;
  wire [8:0] _T_38;
  wire [7:0] _T_40;
  wire [32:0] _T_42;
  wire [31:0] _T_43;
  wire [8:0] _T_44;
  wire [7:0] _T_46;
  wire  _GEN_22;
  wire  _GEN_26;
  wire  _GEN_32;
  wire [8:0] _T_48;
  wire [7:0] _GEN_43;
  wire [8:0] _T_54;
  wire [8:0] _T_56;
  wire [15:0] _T_58;
  wire [15:0] _GEN_48;
  wire [8:0] _T_63;
  wire [8:0] _T_68;
  wire [8:0] _T_73;
  wire [8:0] _T_75;
  wire [15:0] _T_77;
  wire [15:0] _T_78;
  wire [31:0] _T_79;
  wire [31:0] _GEN_55;
  wire  _GEN_58;
  wire  _GEN_62;
  wire  _GEN_66;
  wire  _T_81;
  wire [31:0] _GEN_70;
  assign io_res = _GEN_70;
  assign data_mem__T_49_addr = _T_48;
  assign data_mem__T_49_data = data_mem[data_mem__T_49_addr];
  assign data_mem__T_55_addr = _T_54;
  assign data_mem__T_55_data = data_mem[data_mem__T_55_addr];
  assign data_mem__T_57_addr = _T_56;
  assign data_mem__T_57_data = data_mem[data_mem__T_57_addr];
  assign data_mem__T_64_addr = _T_63;
  assign data_mem__T_64_data = data_mem[data_mem__T_64_addr];
  assign data_mem__T_69_addr = _T_68;
  assign data_mem__T_69_data = data_mem[data_mem__T_69_addr];
  assign data_mem__T_74_addr = _T_73;
  assign data_mem__T_74_data = data_mem[data_mem__T_74_addr];
  assign data_mem__T_76_addr = _T_75;
  assign data_mem__T_76_data = data_mem[data_mem__T_76_addr];
  assign data_mem__T_13_data = _T_14;
  assign data_mem__T_13_addr = _T_12;
  assign data_mem__T_13_mask = _GEN_22;
  assign data_mem__T_13_en = _GEN_22;
  assign data_mem__T_17_data = _T_18;
  assign data_mem__T_17_addr = _T_16;
  assign data_mem__T_17_mask = _GEN_26;
  assign data_mem__T_17_en = _GEN_26;
  assign data_mem__T_23_data = _T_24;
  assign data_mem__T_23_addr = _T_22;
  assign data_mem__T_23_mask = _GEN_26;
  assign data_mem__T_23_en = _GEN_26;
  assign data_mem__T_27_data = _T_28;
  assign data_mem__T_27_addr = _T_26;
  assign data_mem__T_27_mask = _GEN_32;
  assign data_mem__T_27_en = _GEN_32;
  assign data_mem__T_33_data = _T_34;
  assign data_mem__T_33_addr = _T_32;
  assign data_mem__T_33_mask = _GEN_32;
  assign data_mem__T_33_en = _GEN_32;
  assign data_mem__T_39_data = _T_40;
  assign data_mem__T_39_addr = _T_38;
  assign data_mem__T_39_mask = _GEN_32;
  assign data_mem__T_39_en = _GEN_32;
  assign data_mem__T_45_data = _T_46;
  assign data_mem__T_45_addr = _T_44;
  assign data_mem__T_45_mask = _GEN_32;
  assign data_mem__T_45_en = _GEN_32;
  assign _T_11 = 3'h0 == io_mem_func;
  assign _T_12 = io_op_op1[8:0];
  assign _T_14 = io_op_op2[7:0];
  assign _T_15 = 3'h1 == io_mem_func;
  assign _T_16 = io_op_op1[8:0];
  assign _T_18 = io_op_op2[7:0];
  assign _T_20 = io_op_op1 + 32'h1;
  assign _T_21 = _T_20[31:0];
  assign _T_22 = _T_21[8:0];
  assign _T_24 = io_op_op2[15:8];
  assign _T_25 = 3'h2 == io_mem_func;
  assign _T_26 = io_op_op1[8:0];
  assign _T_28 = io_op_op2[7:0];
  assign _T_32 = _T_21[8:0];
  assign _T_34 = io_op_op2[15:8];
  assign _T_36 = io_op_op1 + 32'h2;
  assign _T_37 = _T_36[31:0];
  assign _T_38 = _T_37[8:0];
  assign _T_40 = io_op_op2[23:16];
  assign _T_42 = io_op_op1 + 32'h3;
  assign _T_43 = _T_42[31:0];
  assign _T_44 = _T_43[8:0];
  assign _T_46 = io_op_op2[31:24];
  assign _GEN_22 = io_mem_write ? _T_11 : 1'h0;
  assign _GEN_26 = io_mem_write ? _T_15 : 1'h0;
  assign _GEN_32 = io_mem_write ? _T_25 : 1'h0;
  assign _T_48 = io_op_op1[8:0];
  assign _GEN_43 = data_mem__T_49_data;
  assign _T_54 = _T_21[8:0];
  assign _T_56 = io_op_op1[8:0];
  assign _T_58 = {data_mem__T_55_data,data_mem__T_57_data};
  assign _GEN_48 = _T_15 ? _T_58 : {{8'd0}, _GEN_43};
  assign _T_63 = _T_43[8:0];
  assign _T_68 = _T_37[8:0];
  assign _T_73 = _T_21[8:0];
  assign _T_75 = io_op_op1[8:0];
  assign _T_77 = {data_mem__T_74_data,data_mem__T_76_data};
  assign _T_78 = {data_mem__T_64_data,data_mem__T_69_data};
  assign _T_79 = {_T_78,_T_77};
  assign _GEN_55 = _T_25 ? _T_79 : {{16'd0}, _GEN_48};
  assign _GEN_58 = io_mem_read ? _T_11 : 1'h0;
  assign _GEN_62 = io_mem_read ? _T_15 : 1'h0;
  assign _GEN_66 = io_mem_read ? _T_25 : 1'h0;
  assign _T_81 = io_mem_read == 1'h0;
  assign _GEN_70 = _T_81 ? 32'h0 : _GEN_55;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_mem[initvar] = _GEN_0[7:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if(data_mem__T_13_en & data_mem__T_13_mask) begin
      data_mem[data_mem__T_13_addr] <= data_mem__T_13_data;
    end
    if(data_mem__T_17_en & data_mem__T_17_mask) begin
      data_mem[data_mem__T_17_addr] <= data_mem__T_17_data;
    end
    if(data_mem__T_23_en & data_mem__T_23_mask) begin
      data_mem[data_mem__T_23_addr] <= data_mem__T_23_data;
    end
    if(data_mem__T_27_en & data_mem__T_27_mask) begin
      data_mem[data_mem__T_27_addr] <= data_mem__T_27_data;
    end
    if(data_mem__T_33_en & data_mem__T_33_mask) begin
      data_mem[data_mem__T_33_addr] <= data_mem__T_33_data;
    end
    if(data_mem__T_39_en & data_mem__T_39_mask) begin
      data_mem[data_mem__T_39_addr] <= data_mem__T_39_data;
    end
    if(data_mem__T_45_en & data_mem__T_45_mask) begin
      data_mem[data_mem__T_45_addr] <= data_mem__T_45_data;
    end
  end
endmodule
module ForwardingUnit(
  input        io_reg_w_mem,
  input        io_reg_w_wb,
  input  [4:0] io_rs_rs1,
  input  [4:0] io_rs_rs2,
  input  [4:0] io_rd_mem,
  input  [4:0] io_rd_wb,
  output [1:0] io_fwd_rs1,
  output [1:0] io_fwd_rs2
);
  wire  _T_10;
  wire  _T_11;
  wire  _T_12;
  wire  _T_13;
  wire  _T_14;
  wire  _T_15;
  wire  _T_16;
  wire  _T_17;
  wire  _T_19;
  wire  _T_20;
  wire [1:0] _GEN_1;
  wire  _T_24;
  wire  _T_25;
  wire [1:0] _GEN_2;
  wire  _T_28;
  wire  _T_29;
  wire  _T_32;
  wire  _T_33;
  wire  _T_35;
  wire  _T_36;
  wire [1:0] _GEN_4;
  wire  _T_40;
  wire  _T_41;
  wire [1:0] _GEN_5;
  assign io_fwd_rs1 = _GEN_2;
  assign io_fwd_rs2 = _GEN_5;
  assign _T_10 = io_rd_mem != 5'h0;
  assign _T_11 = io_reg_w_mem & _T_10;
  assign _T_12 = io_rd_mem == io_rs_rs1;
  assign _T_13 = _T_11 & _T_12;
  assign _T_14 = io_rd_wb != 5'h0;
  assign _T_15 = io_reg_w_wb & _T_14;
  assign _T_16 = io_rd_wb == io_rs_rs1;
  assign _T_17 = _T_15 & _T_16;
  assign _T_19 = _T_13 == 1'h0;
  assign _T_20 = _T_19 & _T_17;
  assign _GEN_1 = _T_20 ? 2'h1 : 2'h2;
  assign _T_24 = _T_17 == 1'h0;
  assign _T_25 = _T_19 & _T_24;
  assign _GEN_2 = _T_25 ? 2'h0 : _GEN_1;
  assign _T_28 = io_rd_mem == io_rs_rs2;
  assign _T_29 = _T_11 & _T_28;
  assign _T_32 = io_rd_wb == io_rs_rs2;
  assign _T_33 = _T_15 & _T_32;
  assign _T_35 = _T_29 == 1'h0;
  assign _T_36 = _T_35 & _T_33;
  assign _GEN_4 = _T_36 ? 2'h1 : 2'h2;
  assign _T_40 = _T_33 == 1'h0;
  assign _T_41 = _T_35 & _T_40;
  assign _GEN_5 = _T_41 ? 2'h0 : _GEN_4;
endmodule
module Tx(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  output       io_txd
);
  reg [8:0] data;
  reg [31:0] _GEN_13;
  reg [31:0] ticks;
  reg [31:0] _GEN_14;
  reg [3:0] state;
  reg [31:0] _GEN_15;
  wire  _T_15;
  wire  _T_16;
  wire [8:0] _T_18;
  wire [8:0] _GEN_0;
  wire [31:0] _GEN_1;
  wire [3:0] _GEN_2;
  wire [8:0] _GEN_3;
  wire [31:0] _GEN_4;
  wire [3:0] _GEN_5;
  wire  _T_19;
  wire  _T_20;
  wire  _T_21;
  wire  _T_22;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_26;
  wire  _T_27;
  wire  _T_28;
  wire  _T_29;
  wire  _T_30;
  wire  _T_31;
  wire  _T_32;
  wire  _T_33;
  wire  _T_34;
  wire  _T_35;
  wire  _T_36;
  wire  _T_37;
  wire  _T_38;
  wire  _T_39;
  wire  _T_40;
  wire [7:0] _T_42;
  wire [8:0] _T_43;
  wire [4:0] _T_45;
  wire [4:0] _T_46;
  wire [3:0] _T_47;
  wire [8:0] _GEN_6;
  wire [31:0] _GEN_7;
  wire [3:0] _GEN_8;
  wire  _T_49;
  wire [32:0] _T_51;
  wire [31:0] _T_52;
  wire [31:0] _GEN_9;
  wire [8:0] _GEN_10;
  wire [31:0] _GEN_11;
  wire [3:0] _GEN_12;
  wire  _T_53;
  assign io_enq_ready = _T_15;
  assign io_txd = _T_53;
  assign _T_15 = state == 4'h0;
  assign _T_16 = 4'h0 == state;
  assign _T_18 = {io_enq_bits,1'h0};
  assign _GEN_0 = io_enq_valid ? _T_18 : data;
  assign _GEN_1 = io_enq_valid ? 32'h0 : ticks;
  assign _GEN_2 = io_enq_valid ? 4'hb : state;
  assign _GEN_3 = _T_16 ? _GEN_0 : data;
  assign _GEN_4 = _T_16 ? _GEN_1 : ticks;
  assign _GEN_5 = _T_16 ? _GEN_2 : state;
  assign _T_19 = 4'h1 == state;
  assign _T_20 = 4'h2 == state;
  assign _T_21 = 4'h3 == state;
  assign _T_22 = 4'h4 == state;
  assign _T_23 = 4'h5 == state;
  assign _T_24 = 4'h6 == state;
  assign _T_25 = 4'h7 == state;
  assign _T_26 = 4'h8 == state;
  assign _T_27 = 4'h9 == state;
  assign _T_28 = 4'ha == state;
  assign _T_29 = 4'hb == state;
  assign _T_30 = _T_19 | _T_20;
  assign _T_31 = _T_30 | _T_21;
  assign _T_32 = _T_31 | _T_22;
  assign _T_33 = _T_32 | _T_23;
  assign _T_34 = _T_33 | _T_24;
  assign _T_35 = _T_34 | _T_25;
  assign _T_36 = _T_35 | _T_26;
  assign _T_37 = _T_36 | _T_27;
  assign _T_38 = _T_37 | _T_28;
  assign _T_39 = _T_38 | _T_29;
  assign _T_40 = ticks == 32'h1b2;
  assign _T_42 = data[8:1];
  assign _T_43 = {1'h1,_T_42};
  assign _T_45 = state - 4'h1;
  assign _T_46 = $unsigned(_T_45);
  assign _T_47 = _T_46[3:0];
  assign _GEN_6 = _T_40 ? _T_43 : _GEN_3;
  assign _GEN_7 = _T_40 ? 32'h0 : _GEN_4;
  assign _GEN_8 = _T_40 ? _T_47 : _GEN_5;
  assign _T_49 = _T_40 == 1'h0;
  assign _T_51 = ticks + 32'h1;
  assign _T_52 = _T_51[31:0];
  assign _GEN_9 = _T_49 ? _T_52 : _GEN_7;
  assign _GEN_10 = _T_39 ? _GEN_6 : _GEN_3;
  assign _GEN_11 = _T_39 ? _GEN_9 : _GEN_4;
  assign _GEN_12 = _T_39 ? _GEN_8 : _GEN_5;
  assign _T_53 = data[0];
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_13 = {1{$random}};
  data = _GEN_13[8:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_14 = {1{$random}};
  ticks = _GEN_14[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_15 = {1{$random}};
  state = _GEN_15[3:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (reset) begin
      data <= 9'h1ff;
    end else begin
      if (_T_39) begin
        if (_T_40) begin
          data <= _T_43;
        end else begin
          if (_T_16) begin
            if (io_enq_valid) begin
              data <= _T_18;
            end
          end
        end
      end else begin
        if (_T_16) begin
          if (io_enq_valid) begin
            data <= _T_18;
          end
        end
      end
    end
    if (reset) begin
      ticks <= 32'h0;
    end else begin
      if (_T_39) begin
        if (_T_49) begin
          ticks <= _T_52;
        end else begin
          if (_T_40) begin
            ticks <= 32'h0;
          end else begin
            if (_T_16) begin
              if (io_enq_valid) begin
                ticks <= 32'h0;
              end
            end
          end
        end
      end else begin
        if (_T_16) begin
          if (io_enq_valid) begin
            ticks <= 32'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 4'h0;
    end else begin
      if (_T_39) begin
        if (_T_40) begin
          state <= _T_47;
        end else begin
          if (_T_16) begin
            if (io_enq_valid) begin
              state <= 4'hb;
            end
          end
        end
      end else begin
        if (_T_16) begin
          if (io_enq_valid) begin
            state <= 4'hb;
          end
        end
      end
    end
  end
endmodule
module UART(
  input        clock,
  input        reset,
  input  [7:0] io_in,
  output       io_valid,
  output       io_txd,
  output [7:0] io_r0,
  output [7:0] io_r1,
  output [7:0] io_r2,
  output [7:0] io_r3
);
  wire  tx_clock;
  wire  tx_reset;
  wire  tx_io_enq_ready;
  wire  tx_io_enq_valid;
  wire [7:0] tx_io_enq_bits;
  wire  tx_io_txd;
  wire [7:0] _T_15_0;
  wire [7:0] _T_15_1;
  wire [7:0] _T_15_2;
  wire [7:0] _T_15_3;
  reg [7:0] q_0;
  reg [31:0] _GEN_14;
  reg [7:0] q_1;
  reg [31:0] _GEN_17;
  reg [7:0] q_2;
  reg [31:0] _GEN_20;
  reg [7:0] q_3;
  reg [31:0] _GEN_21;
  reg [1:0] ptr;
  reg [31:0] _GEN_22;
  reg [1:0] cnt;
  reg [31:0] _GEN_23;
  wire [2:0] _T_53;
  wire [1:0] _T_54;
  reg [3:0] i;
  reg [31:0] _GEN_24;
  wire  _T_74;
  wire [2:0] _GEN_19;
  wire  _T_76;
  wire  _T_77;
  wire [1:0] _T_81;
  wire [7:0] _GEN_0;
  wire [7:0] _GEN_2;
  wire [7:0] _GEN_3;
  wire [7:0] _GEN_4;
  wire [7:0] _GEN_5;
  wire [2:0] _T_83;
  wire [1:0] _T_84;
  wire [7:0] _GEN_6;
  wire [7:0] _GEN_7;
  wire [7:0] _GEN_8;
  wire [7:0] _GEN_9;
  wire [1:0] _GEN_10;
  wire  _T_86;
  wire  _T_87;
  wire [7:0] _GEN_1;
  wire [7:0] _GEN_11;
  wire [7:0] _GEN_12;
  wire [7:0] _GEN_13;
  wire [2:0] _T_92;
  wire [2:0] _T_93;
  wire [1:0] _T_94;
  wire [2:0] _T_96;
  wire [1:0] _T_97;
  wire [1:0] _GEN_15;
  wire [1:0] _GEN_16;
  wire  _T_104;
  wire  _T_105;
  wire  _T_107;
  wire  _GEN_18;
  Tx tx (
    .clock(tx_clock),
    .reset(tx_reset),
    .io_enq_ready(tx_io_enq_ready),
    .io_enq_valid(tx_io_enq_valid),
    .io_enq_bits(tx_io_enq_bits),
    .io_txd(tx_io_txd)
  );
  assign io_valid = _GEN_18;
  assign io_txd = tx_io_txd;
  assign io_r0 = q_0;
  assign io_r1 = q_1;
  assign io_r2 = q_2;
  assign io_r3 = q_3;
  assign tx_clock = clock;
  assign tx_reset = reset;
  assign tx_io_enq_valid = _T_86;
  assign tx_io_enq_bits = _GEN_1;
  assign _T_15_0 = 8'h0;
  assign _T_15_1 = 8'h0;
  assign _T_15_2 = 8'h0;
  assign _T_15_3 = 8'h0;
  assign _T_53 = ptr + cnt;
  assign _T_54 = _T_53[1:0];
  assign _T_74 = io_in != 8'h0;
  assign _GEN_19 = {{1'd0}, cnt};
  assign _T_76 = _GEN_19 != 3'h4;
  assign _T_77 = _T_74 & _T_76;
  assign _T_81 = i[1:0];
  assign _GEN_0 = io_in;
  assign _GEN_2 = 2'h0 == _T_81 ? _GEN_0 : q_0;
  assign _GEN_3 = 2'h1 == _T_81 ? _GEN_0 : q_1;
  assign _GEN_4 = 2'h2 == _T_81 ? _GEN_0 : q_2;
  assign _GEN_5 = 2'h3 == _T_81 ? _GEN_0 : q_3;
  assign _T_83 = cnt + 2'h1;
  assign _T_84 = _T_83[1:0];
  assign _GEN_6 = _T_77 ? _GEN_2 : q_0;
  assign _GEN_7 = _T_77 ? _GEN_3 : q_1;
  assign _GEN_8 = _T_77 ? _GEN_4 : q_2;
  assign _GEN_9 = _T_77 ? _GEN_5 : q_3;
  assign _GEN_10 = _T_77 ? _T_84 : cnt;
  assign _T_86 = cnt != 2'h0;
  assign _T_87 = tx_io_enq_ready & _T_86;
  assign _GEN_1 = _GEN_13;
  assign _GEN_11 = 2'h1 == ptr ? q_1 : q_0;
  assign _GEN_12 = 2'h2 == ptr ? q_2 : _GEN_11;
  assign _GEN_13 = 2'h3 == ptr ? q_3 : _GEN_12;
  assign _T_92 = cnt - 2'h1;
  assign _T_93 = $unsigned(_T_92);
  assign _T_94 = _T_93[1:0];
  assign _T_96 = ptr + 2'h1;
  assign _T_97 = _T_96[1:0];
  assign _GEN_15 = _T_87 ? _T_94 : _GEN_10;
  assign _GEN_16 = _T_87 ? _T_97 : ptr;
  assign _T_104 = _T_74 | _T_86;
  assign _T_105 = _T_104 & tx_io_enq_ready;
  assign _T_107 = _T_105 == 1'h0;
  assign _GEN_18 = _T_107 ? tx_io_enq_ready : 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_14 = {1{$random}};
  q_0 = _GEN_14[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_17 = {1{$random}};
  q_1 = _GEN_17[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_20 = {1{$random}};
  q_2 = _GEN_20[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_21 = {1{$random}};
  q_3 = _GEN_21[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_22 = {1{$random}};
  ptr = _GEN_22[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_23 = {1{$random}};
  cnt = _GEN_23[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_24 = {1{$random}};
  i = _GEN_24[3:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if (reset) begin
      q_0 <= _T_15_0;
    end else begin
      if (_T_77) begin
        if (2'h0 == _T_81) begin
          q_0 <= _GEN_0;
        end
      end
    end
    if (reset) begin
      q_1 <= _T_15_1;
    end else begin
      if (_T_77) begin
        if (2'h1 == _T_81) begin
          q_1 <= _GEN_0;
        end
      end
    end
    if (reset) begin
      q_2 <= _T_15_2;
    end else begin
      if (_T_77) begin
        if (2'h2 == _T_81) begin
          q_2 <= _GEN_0;
        end
      end
    end
    if (reset) begin
      q_3 <= _T_15_3;
    end else begin
      if (_T_77) begin
        if (2'h3 == _T_81) begin
          q_3 <= _GEN_0;
        end
      end
    end
    if (reset) begin
      ptr <= 2'h0;
    end else begin
      if (_T_87) begin
        ptr <= _T_97;
      end
    end
    if (reset) begin
      cnt <= 2'h0;
    end else begin
      if (_T_87) begin
        cnt <= _T_94;
      end else begin
        if (_T_77) begin
          cnt <= _T_84;
        end
      end
    end
    if (reset) begin
      i <= {{2'd0}, _T_54};
    end else begin
      i <= {{2'd0}, _T_54};
    end
  end
endmodule
module PipelineIF_ID(
  input         clock,
  input  [31:0] io_in_pc_next,
  input  [31:0] io_in_inst,
  output [31:0] io_out_pc_next,
  output [31:0] io_out_inst
);
  reg [31:0] _T_12_pc_next;
  reg [31:0] _GEN_0;
  reg [31:0] _T_12_inst;
  reg [31:0] _GEN_1;
  assign io_out_pc_next = _T_12_pc_next;
  assign io_out_inst = _T_12_inst;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_0 = {1{$random}};
  _T_12_pc_next = _GEN_0[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1 = {1{$random}};
  _T_12_inst = _GEN_1[31:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    _T_12_pc_next <= io_in_pc_next;
    _T_12_inst <= io_in_inst;
  end
endmodule
module PipelineID_EX(
  input         clock,
  input         io_in_WB_reg_w,
  input         io_in_WB_rd_mem,
  input         io_in_MEM_write,
  input         io_in_MEM_read,
  input  [2:0]  io_in_MEM_func,
  input  [6:0]  io_in_EX_opcode,
  input         io_in_EX_alu_sel,
  input         io_in_EX_dst_sel,
  input  [2:0]  io_in_EX_alu_op_func,
  input         io_in_EX_alu_op_alt,
  input  [31:0] io_in_op_op1,
  input  [31:0] io_in_op_op2,
  input  [4:0]  io_in_rs_rs1,
  input  [4:0]  io_in_rs_rs2,
  input  [4:0]  io_in_rd,
  input  [31:0] io_in_imm,
  input  [31:0] io_in_pc_next,
  output        io_out_WB_reg_w,
  output        io_out_WB_rd_mem,
  output        io_out_MEM_write,
  output        io_out_MEM_read,
  output [2:0]  io_out_MEM_func,
  output [6:0]  io_out_EX_opcode,
  output        io_out_EX_alu_sel,
  output        io_out_EX_dst_sel,
  output [2:0]  io_out_EX_alu_op_func,
  output        io_out_EX_alu_op_alt,
  output [31:0] io_out_op_op1,
  output [31:0] io_out_op_op2,
  output [4:0]  io_out_rs_rs1,
  output [4:0]  io_out_rs_rs2,
  output [4:0]  io_out_rd,
  output [31:0] io_out_imm,
  output [31:0] io_out_pc_next
);
  reg  _T_76_WB_reg_w;
  reg [31:0] _GEN_0;
  reg  _T_76_WB_rd_mem;
  reg [31:0] _GEN_1;
  reg  _T_76_MEM_write;
  reg [31:0] _GEN_2;
  reg  _T_76_MEM_read;
  reg [31:0] _GEN_3;
  reg [2:0] _T_76_MEM_func;
  reg [31:0] _GEN_4;
  reg [6:0] _T_76_EX_opcode;
  reg [31:0] _GEN_5;
  reg  _T_76_EX_alu_sel;
  reg [31:0] _GEN_6;
  reg  _T_76_EX_dst_sel;
  reg [31:0] _GEN_7;
  reg [2:0] _T_76_EX_alu_op_func;
  reg [31:0] _GEN_8;
  reg  _T_76_EX_alu_op_alt;
  reg [31:0] _GEN_9;
  reg [31:0] _T_76_op_op1;
  reg [31:0] _GEN_10;
  reg [31:0] _T_76_op_op2;
  reg [31:0] _GEN_11;
  reg [4:0] _T_76_rs_rs1;
  reg [31:0] _GEN_12;
  reg [4:0] _T_76_rs_rs2;
  reg [31:0] _GEN_13;
  reg [4:0] _T_76_rd;
  reg [31:0] _GEN_14;
  reg [31:0] _T_76_imm;
  reg [31:0] _GEN_15;
  reg [31:0] _T_76_pc_next;
  reg [31:0] _GEN_16;
  assign io_out_WB_reg_w = _T_76_WB_reg_w;
  assign io_out_WB_rd_mem = _T_76_WB_rd_mem;
  assign io_out_MEM_write = _T_76_MEM_write;
  assign io_out_MEM_read = _T_76_MEM_read;
  assign io_out_MEM_func = _T_76_MEM_func;
  assign io_out_EX_opcode = _T_76_EX_opcode;
  assign io_out_EX_alu_sel = _T_76_EX_alu_sel;
  assign io_out_EX_dst_sel = _T_76_EX_dst_sel;
  assign io_out_EX_alu_op_func = _T_76_EX_alu_op_func;
  assign io_out_EX_alu_op_alt = _T_76_EX_alu_op_alt;
  assign io_out_op_op1 = _T_76_op_op1;
  assign io_out_op_op2 = _T_76_op_op2;
  assign io_out_rs_rs1 = _T_76_rs_rs1;
  assign io_out_rs_rs2 = _T_76_rs_rs2;
  assign io_out_rd = _T_76_rd;
  assign io_out_imm = _T_76_imm;
  assign io_out_pc_next = _T_76_pc_next;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_0 = {1{$random}};
  _T_76_WB_reg_w = _GEN_0[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1 = {1{$random}};
  _T_76_WB_rd_mem = _GEN_1[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2 = {1{$random}};
  _T_76_MEM_write = _GEN_2[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_3 = {1{$random}};
  _T_76_MEM_read = _GEN_3[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_4 = {1{$random}};
  _T_76_MEM_func = _GEN_4[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_5 = {1{$random}};
  _T_76_EX_opcode = _GEN_5[6:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_6 = {1{$random}};
  _T_76_EX_alu_sel = _GEN_6[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_7 = {1{$random}};
  _T_76_EX_dst_sel = _GEN_7[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_8 = {1{$random}};
  _T_76_EX_alu_op_func = _GEN_8[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_9 = {1{$random}};
  _T_76_EX_alu_op_alt = _GEN_9[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_10 = {1{$random}};
  _T_76_op_op1 = _GEN_10[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_11 = {1{$random}};
  _T_76_op_op2 = _GEN_11[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_12 = {1{$random}};
  _T_76_rs_rs1 = _GEN_12[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_13 = {1{$random}};
  _T_76_rs_rs2 = _GEN_13[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_14 = {1{$random}};
  _T_76_rd = _GEN_14[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_15 = {1{$random}};
  _T_76_imm = _GEN_15[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_16 = {1{$random}};
  _T_76_pc_next = _GEN_16[31:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    _T_76_WB_reg_w <= io_in_WB_reg_w;
    _T_76_WB_rd_mem <= io_in_WB_rd_mem;
    _T_76_MEM_write <= io_in_MEM_write;
    _T_76_MEM_read <= io_in_MEM_read;
    _T_76_MEM_func <= io_in_MEM_func;
    _T_76_EX_opcode <= io_in_EX_opcode;
    _T_76_EX_alu_sel <= io_in_EX_alu_sel;
    _T_76_EX_dst_sel <= io_in_EX_dst_sel;
    _T_76_EX_alu_op_func <= io_in_EX_alu_op_func;
    _T_76_EX_alu_op_alt <= io_in_EX_alu_op_alt;
    _T_76_op_op1 <= io_in_op_op1;
    _T_76_op_op2 <= io_in_op_op2;
    _T_76_rs_rs1 <= io_in_rs_rs1;
    _T_76_rs_rs2 <= io_in_rs_rs2;
    _T_76_rd <= io_in_rd;
    _T_76_imm <= io_in_imm;
    _T_76_pc_next <= io_in_pc_next;
  end
endmodule
module PipelineEX_MEM(
  input         clock,
  input         io_in_WB_reg_w,
  input         io_in_WB_rd_mem,
  input         io_in_MEM_write,
  input         io_in_MEM_read,
  input  [2:0]  io_in_MEM_func,
  input  [31:0] io_in_op_op1,
  input  [31:0] io_in_op_op2,
  input  [4:0]  io_in_rd,
  input  [31:0] io_in_pc_next,
  output        io_out_WB_reg_w,
  output        io_out_WB_rd_mem,
  output        io_out_MEM_write,
  output        io_out_MEM_read,
  output [2:0]  io_out_MEM_func,
  output [31:0] io_out_op_op1,
  output [31:0] io_out_op_op2,
  output [4:0]  io_out_rd,
  output [31:0] io_out_pc_next
);
  reg  _T_48_WB_reg_w;
  reg [31:0] _GEN_0;
  reg  _T_48_WB_rd_mem;
  reg [31:0] _GEN_1;
  reg  _T_48_MEM_write;
  reg [31:0] _GEN_2;
  reg  _T_48_MEM_read;
  reg [31:0] _GEN_3;
  reg [2:0] _T_48_MEM_func;
  reg [31:0] _GEN_4;
  reg [31:0] _T_48_op_op1;
  reg [31:0] _GEN_5;
  reg [31:0] _T_48_op_op2;
  reg [31:0] _GEN_6;
  reg [4:0] _T_48_rd;
  reg [31:0] _GEN_7;
  reg [31:0] _T_48_pc_next;
  reg [31:0] _GEN_8;
  assign io_out_WB_reg_w = _T_48_WB_reg_w;
  assign io_out_WB_rd_mem = _T_48_WB_rd_mem;
  assign io_out_MEM_write = _T_48_MEM_write;
  assign io_out_MEM_read = _T_48_MEM_read;
  assign io_out_MEM_func = _T_48_MEM_func;
  assign io_out_op_op1 = _T_48_op_op1;
  assign io_out_op_op2 = _T_48_op_op2;
  assign io_out_rd = _T_48_rd;
  assign io_out_pc_next = _T_48_pc_next;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_0 = {1{$random}};
  _T_48_WB_reg_w = _GEN_0[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1 = {1{$random}};
  _T_48_WB_rd_mem = _GEN_1[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2 = {1{$random}};
  _T_48_MEM_write = _GEN_2[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_3 = {1{$random}};
  _T_48_MEM_read = _GEN_3[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_4 = {1{$random}};
  _T_48_MEM_func = _GEN_4[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_5 = {1{$random}};
  _T_48_op_op1 = _GEN_5[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_6 = {1{$random}};
  _T_48_op_op2 = _GEN_6[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_7 = {1{$random}};
  _T_48_rd = _GEN_7[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_8 = {1{$random}};
  _T_48_pc_next = _GEN_8[31:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    _T_48_WB_reg_w <= io_in_WB_reg_w;
    _T_48_WB_rd_mem <= io_in_WB_rd_mem;
    _T_48_MEM_write <= io_in_MEM_write;
    _T_48_MEM_read <= io_in_MEM_read;
    _T_48_MEM_func <= io_in_MEM_func;
    _T_48_op_op1 <= io_in_op_op1;
    _T_48_op_op2 <= io_in_op_op2;
    _T_48_rd <= io_in_rd;
    _T_48_pc_next <= io_in_pc_next;
  end
endmodule
module PipelineMEM_WB(
  input         clock,
  input         io_in_WB_reg_w,
  input         io_in_WB_rd_mem,
  input  [31:0] io_in_alu_res,
  input  [31:0] io_in_mem_res,
  input  [4:0]  io_in_rd,
  output        io_out_WB_reg_w,
  output        io_out_WB_rd_mem,
  output [31:0] io_out_alu_res,
  output [31:0] io_out_mem_res,
  output [4:0]  io_out_rd
);
  reg  _T_24_WB_reg_w;
  reg [31:0] _GEN_0;
  reg  _T_24_WB_rd_mem;
  reg [31:0] _GEN_1;
  reg [31:0] _T_24_alu_res;
  reg [31:0] _GEN_2;
  reg [31:0] _T_24_mem_res;
  reg [31:0] _GEN_3;
  reg [4:0] _T_24_rd;
  reg [31:0] _GEN_4;
  assign io_out_WB_reg_w = _T_24_WB_reg_w;
  assign io_out_WB_rd_mem = _T_24_WB_rd_mem;
  assign io_out_alu_res = _T_24_alu_res;
  assign io_out_mem_res = _T_24_mem_res;
  assign io_out_rd = _T_24_rd;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_0 = {1{$random}};
  _T_24_WB_reg_w = _GEN_0[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_1 = {1{$random}};
  _T_24_WB_rd_mem = _GEN_1[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_2 = {1{$random}};
  _T_24_alu_res = _GEN_2[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_3 = {1{$random}};
  _T_24_mem_res = _GEN_3[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_4 = {1{$random}};
  _T_24_rd = _GEN_4[4:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    _T_24_WB_reg_w <= io_in_WB_reg_w;
    _T_24_WB_rd_mem <= io_in_WB_rd_mem;
    _T_24_alu_res <= io_in_alu_res;
    _T_24_mem_res <= io_in_mem_res;
    _T_24_rd <= io_in_rd;
  end
endmodule
module CPU(
  input         clock,
  input         reset,
  output        io_txd,
  output [7:0]  io_r0,
  output [7:0]  io_r1,
  output [7:0]  io_r2,
  output [7:0]  io_r3,
  output [31:0] io_inst
);
  wire  instMem_clock;
  wire [31:0] instMem_io_pc;
  wire [31:0] instMem_io_inst;
  wire  counter_clock;
  wire  counter_reset;
  wire  counter_io_branch;
  wire [31:0] counter_io_pc_src;
  wire [31:0] counter_io_pc_next;
  wire [31:0] counter_io_pc;
  wire [31:0] decoder_io_inst;
  wire [6:0] decoder_io_ctrl_opcode;
  wire [2:0] decoder_io_ctrl_funct3;
  wire [6:0] decoder_io_ctrl_funct7;
  wire [4:0] decoder_io_rs_rs1;
  wire [4:0] decoder_io_rs_rs2;
  wire [4:0] decoder_io_rd;
  wire [31:0] decoder_io_imm;
  wire [6:0] control_io_ctrl_opcode;
  wire [2:0] control_io_ctrl_funct3;
  wire [6:0] control_io_ctrl_funct7;
  wire  control_io_WB_reg_w;
  wire  control_io_WB_rd_mem;
  wire  control_io_MEM_branch;
  wire  control_io_MEM_write;
  wire  control_io_MEM_read;
  wire [2:0] control_io_MEM_func;
  wire [6:0] control_io_EX_opcode;
  wire  control_io_EX_alu_sel;
  wire  control_io_EX_dst_sel;
  wire [2:0] control_io_EX_alu_op_func;
  wire  control_io_EX_alu_op_alt;
  wire  regs_clock;
  wire [4:0] regs_io_rs_rs1;
  wire [4:0] regs_io_rs_rs2;
  wire  regs_io_reg_w;
  wire [4:0] regs_io_rd;
  wire [31:0] regs_io_res;
  wire [31:0] regs_io_op_op1;
  wire [31:0] regs_io_op_op2;
  wire [6:0] alu_io_opcode;
  wire [2:0] alu_io_alu_op_func;
  wire  alu_io_alu_op_alt;
  wire [31:0] alu_io_op_op1;
  wire [31:0] alu_io_op_op2;
  wire [31:0] alu_io_res;
  wire  dataMem_clock;
  wire  dataMem_io_mem_write;
  wire  dataMem_io_mem_read;
  wire [2:0] dataMem_io_mem_func;
  wire [31:0] dataMem_io_op_op1;
  wire [31:0] dataMem_io_op_op2;
  wire [31:0] dataMem_io_res;
  wire  fwdUnit_io_reg_w_mem;
  wire  fwdUnit_io_reg_w_wb;
  wire [4:0] fwdUnit_io_rs_rs1;
  wire [4:0] fwdUnit_io_rs_rs2;
  wire [4:0] fwdUnit_io_rd_mem;
  wire [4:0] fwdUnit_io_rd_wb;
  wire [1:0] fwdUnit_io_fwd_rs1;
  wire [1:0] fwdUnit_io_fwd_rs2;
  wire  uart_clock;
  wire  uart_reset;
  wire [7:0] uart_io_in;
  wire  uart_io_valid;
  wire  uart_io_txd;
  wire [7:0] uart_io_r0;
  wire [7:0] uart_io_r1;
  wire [7:0] uart_io_r2;
  wire [7:0] uart_io_r3;
  wire  IF_ID_clock;
  wire [31:0] IF_ID_io_in_pc_next;
  wire [31:0] IF_ID_io_in_inst;
  wire [31:0] IF_ID_io_out_pc_next;
  wire [31:0] IF_ID_io_out_inst;
  wire  ID_EX_clock;
  wire  ID_EX_io_in_WB_reg_w;
  wire  ID_EX_io_in_WB_rd_mem;
  wire  ID_EX_io_in_MEM_write;
  wire  ID_EX_io_in_MEM_read;
  wire [2:0] ID_EX_io_in_MEM_func;
  wire [6:0] ID_EX_io_in_EX_opcode;
  wire  ID_EX_io_in_EX_alu_sel;
  wire  ID_EX_io_in_EX_dst_sel;
  wire [2:0] ID_EX_io_in_EX_alu_op_func;
  wire  ID_EX_io_in_EX_alu_op_alt;
  wire [31:0] ID_EX_io_in_op_op1;
  wire [31:0] ID_EX_io_in_op_op2;
  wire [4:0] ID_EX_io_in_rs_rs1;
  wire [4:0] ID_EX_io_in_rs_rs2;
  wire [4:0] ID_EX_io_in_rd;
  wire [31:0] ID_EX_io_in_imm;
  wire [31:0] ID_EX_io_in_pc_next;
  wire  ID_EX_io_out_WB_reg_w;
  wire  ID_EX_io_out_WB_rd_mem;
  wire  ID_EX_io_out_MEM_write;
  wire  ID_EX_io_out_MEM_read;
  wire [2:0] ID_EX_io_out_MEM_func;
  wire [6:0] ID_EX_io_out_EX_opcode;
  wire  ID_EX_io_out_EX_alu_sel;
  wire  ID_EX_io_out_EX_dst_sel;
  wire [2:0] ID_EX_io_out_EX_alu_op_func;
  wire  ID_EX_io_out_EX_alu_op_alt;
  wire [31:0] ID_EX_io_out_op_op1;
  wire [31:0] ID_EX_io_out_op_op2;
  wire [4:0] ID_EX_io_out_rs_rs1;
  wire [4:0] ID_EX_io_out_rs_rs2;
  wire [4:0] ID_EX_io_out_rd;
  wire [31:0] ID_EX_io_out_imm;
  wire [31:0] ID_EX_io_out_pc_next;
  wire  EX_MEM_clock;
  wire  EX_MEM_io_in_WB_reg_w;
  wire  EX_MEM_io_in_WB_rd_mem;
  wire  EX_MEM_io_in_MEM_write;
  wire  EX_MEM_io_in_MEM_read;
  wire [2:0] EX_MEM_io_in_MEM_func;
  wire [31:0] EX_MEM_io_in_op_op1;
  wire [31:0] EX_MEM_io_in_op_op2;
  wire [4:0] EX_MEM_io_in_rd;
  wire [31:0] EX_MEM_io_in_pc_next;
  wire  EX_MEM_io_out_WB_reg_w;
  wire  EX_MEM_io_out_WB_rd_mem;
  wire  EX_MEM_io_out_MEM_write;
  wire  EX_MEM_io_out_MEM_read;
  wire [2:0] EX_MEM_io_out_MEM_func;
  wire [31:0] EX_MEM_io_out_op_op1;
  wire [31:0] EX_MEM_io_out_op_op2;
  wire [4:0] EX_MEM_io_out_rd;
  wire [31:0] EX_MEM_io_out_pc_next;
  wire  MEM_WB_clock;
  wire  MEM_WB_io_in_WB_reg_w;
  wire  MEM_WB_io_in_WB_rd_mem;
  wire [31:0] MEM_WB_io_in_alu_res;
  wire [31:0] MEM_WB_io_in_mem_res;
  wire [4:0] MEM_WB_io_in_rd;
  wire  MEM_WB_io_out_WB_reg_w;
  wire  MEM_WB_io_out_WB_rd_mem;
  wire [31:0] MEM_WB_io_out_alu_res;
  wire [31:0] MEM_WB_io_out_mem_res;
  wire [4:0] MEM_WB_io_out_rd;
  wire  _T_51;
  wire  _T_52;
  wire  _T_54;
  wire  _T_55;
  wire [32:0] _T_56;
  wire [31:0] _T_57;
  wire [32:0] _T_59;
  wire [32:0] _T_60;
  wire [31:0] _T_61;
  wire [31:0] _T_62;
  wire [6:0] _T_63;
  wire [2:0] _T_64;
  wire [6:0] _T_65;
  wire  _T_66;
  wire [31:0] _T_67;
  wire  _T_68;
  wire [31:0] _T_69;
  wire  _T_70;
  wire [31:0] _T_71;
  wire [31:0] _T_72;
  wire [31:0] _T_73;
  wire [31:0] _T_74;
  wire  _T_75;
  wire [31:0] _T_76;
  wire  _T_77;
  wire [31:0] _T_78;
  wire  _T_79;
  wire [31:0] _T_80;
  wire [4:0] _T_81;
  wire [31:0] _T_82;
  wire  _T_84;
  wire  _T_85;
  wire [31:0] _GEN_0;
  wire  _T_87;
  wire [31:0] _GEN_1;
  reg [4:0] _GEN_2;
  reg [31:0] _GEN_6;
  reg [4:0] _GEN_3;
  reg [31:0] _GEN_7;
  reg [4:0] _GEN_4;
  reg [31:0] _GEN_8;
  reg  _GEN_5;
  reg [31:0] _GEN_9;
  InstructionMemory instMem (
    .clock(instMem_clock),
    .io_pc(instMem_io_pc),
    .io_inst(instMem_io_inst)
  );
  ProgramCounter counter (
    .clock(counter_clock),
    .reset(counter_reset),
    .io_branch(counter_io_branch),
    .io_pc_src(counter_io_pc_src),
    .io_pc_next(counter_io_pc_next),
    .io_pc(counter_io_pc)
  );
  Decoder decoder (
    .io_inst(decoder_io_inst),
    .io_ctrl_opcode(decoder_io_ctrl_opcode),
    .io_ctrl_funct3(decoder_io_ctrl_funct3),
    .io_ctrl_funct7(decoder_io_ctrl_funct7),
    .io_rs_rs1(decoder_io_rs_rs1),
    .io_rs_rs2(decoder_io_rs_rs2),
    .io_rd(decoder_io_rd),
    .io_imm(decoder_io_imm)
  );
  Control control (
    .io_ctrl_opcode(control_io_ctrl_opcode),
    .io_ctrl_funct3(control_io_ctrl_funct3),
    .io_ctrl_funct7(control_io_ctrl_funct7),
    .io_WB_reg_w(control_io_WB_reg_w),
    .io_WB_rd_mem(control_io_WB_rd_mem),
    .io_MEM_branch(control_io_MEM_branch),
    .io_MEM_write(control_io_MEM_write),
    .io_MEM_read(control_io_MEM_read),
    .io_MEM_func(control_io_MEM_func),
    .io_EX_opcode(control_io_EX_opcode),
    .io_EX_alu_sel(control_io_EX_alu_sel),
    .io_EX_dst_sel(control_io_EX_dst_sel),
    .io_EX_alu_op_func(control_io_EX_alu_op_func),
    .io_EX_alu_op_alt(control_io_EX_alu_op_alt)
  );
  Registers regs (
    .clock(regs_clock),
    .io_rs_rs1(regs_io_rs_rs1),
    .io_rs_rs2(regs_io_rs_rs2),
    .io_reg_w(regs_io_reg_w),
    .io_rd(regs_io_rd),
    .io_res(regs_io_res),
    .io_op_op1(regs_io_op_op1),
    .io_op_op2(regs_io_op_op2)
  );
  ALU alu (
    .io_opcode(alu_io_opcode),
    .io_alu_op_func(alu_io_alu_op_func),
    .io_alu_op_alt(alu_io_alu_op_alt),
    .io_op_op1(alu_io_op_op1),
    .io_op_op2(alu_io_op_op2),
    .io_res(alu_io_res)
  );
  DataMemory dataMem (
    .clock(dataMem_clock),
    .io_mem_write(dataMem_io_mem_write),
    .io_mem_read(dataMem_io_mem_read),
    .io_mem_func(dataMem_io_mem_func),
    .io_op_op1(dataMem_io_op_op1),
    .io_op_op2(dataMem_io_op_op2),
    .io_res(dataMem_io_res)
  );
  ForwardingUnit fwdUnit (
    .io_reg_w_mem(fwdUnit_io_reg_w_mem),
    .io_reg_w_wb(fwdUnit_io_reg_w_wb),
    .io_rs_rs1(fwdUnit_io_rs_rs1),
    .io_rs_rs2(fwdUnit_io_rs_rs2),
    .io_rd_mem(fwdUnit_io_rd_mem),
    .io_rd_wb(fwdUnit_io_rd_wb),
    .io_fwd_rs1(fwdUnit_io_fwd_rs1),
    .io_fwd_rs2(fwdUnit_io_fwd_rs2)
  );
  UART uart (
    .clock(uart_clock),
    .reset(uart_reset),
    .io_in(uart_io_in),
    .io_valid(uart_io_valid),
    .io_txd(uart_io_txd),
    .io_r0(uart_io_r0),
    .io_r1(uart_io_r1),
    .io_r2(uart_io_r2),
    .io_r3(uart_io_r3)
  );
  PipelineIF_ID IF_ID (
    .clock(IF_ID_clock),
    .io_in_pc_next(IF_ID_io_in_pc_next),
    .io_in_inst(IF_ID_io_in_inst),
    .io_out_pc_next(IF_ID_io_out_pc_next),
    .io_out_inst(IF_ID_io_out_inst)
  );
  PipelineID_EX ID_EX (
    .clock(ID_EX_clock),
    .io_in_WB_reg_w(ID_EX_io_in_WB_reg_w),
    .io_in_WB_rd_mem(ID_EX_io_in_WB_rd_mem),
    .io_in_MEM_write(ID_EX_io_in_MEM_write),
    .io_in_MEM_read(ID_EX_io_in_MEM_read),
    .io_in_MEM_func(ID_EX_io_in_MEM_func),
    .io_in_EX_opcode(ID_EX_io_in_EX_opcode),
    .io_in_EX_alu_sel(ID_EX_io_in_EX_alu_sel),
    .io_in_EX_dst_sel(ID_EX_io_in_EX_dst_sel),
    .io_in_EX_alu_op_func(ID_EX_io_in_EX_alu_op_func),
    .io_in_EX_alu_op_alt(ID_EX_io_in_EX_alu_op_alt),
    .io_in_op_op1(ID_EX_io_in_op_op1),
    .io_in_op_op2(ID_EX_io_in_op_op2),
    .io_in_rs_rs1(ID_EX_io_in_rs_rs1),
    .io_in_rs_rs2(ID_EX_io_in_rs_rs2),
    .io_in_rd(ID_EX_io_in_rd),
    .io_in_imm(ID_EX_io_in_imm),
    .io_in_pc_next(ID_EX_io_in_pc_next),
    .io_out_WB_reg_w(ID_EX_io_out_WB_reg_w),
    .io_out_WB_rd_mem(ID_EX_io_out_WB_rd_mem),
    .io_out_MEM_write(ID_EX_io_out_MEM_write),
    .io_out_MEM_read(ID_EX_io_out_MEM_read),
    .io_out_MEM_func(ID_EX_io_out_MEM_func),
    .io_out_EX_opcode(ID_EX_io_out_EX_opcode),
    .io_out_EX_alu_sel(ID_EX_io_out_EX_alu_sel),
    .io_out_EX_dst_sel(ID_EX_io_out_EX_dst_sel),
    .io_out_EX_alu_op_func(ID_EX_io_out_EX_alu_op_func),
    .io_out_EX_alu_op_alt(ID_EX_io_out_EX_alu_op_alt),
    .io_out_op_op1(ID_EX_io_out_op_op1),
    .io_out_op_op2(ID_EX_io_out_op_op2),
    .io_out_rs_rs1(ID_EX_io_out_rs_rs1),
    .io_out_rs_rs2(ID_EX_io_out_rs_rs2),
    .io_out_rd(ID_EX_io_out_rd),
    .io_out_imm(ID_EX_io_out_imm),
    .io_out_pc_next(ID_EX_io_out_pc_next)
  );
  PipelineEX_MEM EX_MEM (
    .clock(EX_MEM_clock),
    .io_in_WB_reg_w(EX_MEM_io_in_WB_reg_w),
    .io_in_WB_rd_mem(EX_MEM_io_in_WB_rd_mem),
    .io_in_MEM_write(EX_MEM_io_in_MEM_write),
    .io_in_MEM_read(EX_MEM_io_in_MEM_read),
    .io_in_MEM_func(EX_MEM_io_in_MEM_func),
    .io_in_op_op1(EX_MEM_io_in_op_op1),
    .io_in_op_op2(EX_MEM_io_in_op_op2),
    .io_in_rd(EX_MEM_io_in_rd),
    .io_in_pc_next(EX_MEM_io_in_pc_next),
    .io_out_WB_reg_w(EX_MEM_io_out_WB_reg_w),
    .io_out_WB_rd_mem(EX_MEM_io_out_WB_rd_mem),
    .io_out_MEM_write(EX_MEM_io_out_MEM_write),
    .io_out_MEM_read(EX_MEM_io_out_MEM_read),
    .io_out_MEM_func(EX_MEM_io_out_MEM_func),
    .io_out_op_op1(EX_MEM_io_out_op_op1),
    .io_out_op_op2(EX_MEM_io_out_op_op2),
    .io_out_rd(EX_MEM_io_out_rd),
    .io_out_pc_next(EX_MEM_io_out_pc_next)
  );
  PipelineMEM_WB MEM_WB (
    .clock(MEM_WB_clock),
    .io_in_WB_reg_w(MEM_WB_io_in_WB_reg_w),
    .io_in_WB_rd_mem(MEM_WB_io_in_WB_rd_mem),
    .io_in_alu_res(MEM_WB_io_in_alu_res),
    .io_in_mem_res(MEM_WB_io_in_mem_res),
    .io_in_rd(MEM_WB_io_in_rd),
    .io_out_WB_reg_w(MEM_WB_io_out_WB_reg_w),
    .io_out_WB_rd_mem(MEM_WB_io_out_WB_rd_mem),
    .io_out_alu_res(MEM_WB_io_out_alu_res),
    .io_out_mem_res(MEM_WB_io_out_mem_res),
    .io_out_rd(MEM_WB_io_out_rd)
  );
  assign io_txd = uart_io_txd;
  assign io_r0 = uart_io_r0;
  assign io_r1 = uart_io_r1;
  assign io_r2 = uart_io_r2;
  assign io_r3 = uart_io_r3;
  assign io_inst = instMem_io_inst;
  assign instMem_clock = clock;
  assign instMem_io_pc = counter_io_pc;
  assign counter_clock = clock;
  assign counter_reset = reset;
  assign counter_io_branch = _T_55;
  assign counter_io_pc_src = _T_62;
  assign decoder_io_inst = IF_ID_io_out_inst;
  assign control_io_ctrl_opcode = _T_63;
  assign control_io_ctrl_funct3 = _T_64;
  assign control_io_ctrl_funct7 = _T_65;
  assign regs_clock = clock;
  assign regs_io_rs_rs1 = decoder_io_rs_rs1;
  assign regs_io_rs_rs2 = decoder_io_rs_rs2;
  assign regs_io_reg_w = MEM_WB_io_out_WB_reg_w;
  assign regs_io_rd = MEM_WB_io_out_rd;
  assign regs_io_res = _T_82;
  assign alu_io_opcode = ID_EX_io_out_EX_opcode;
  assign alu_io_alu_op_func = ID_EX_io_out_EX_alu_op_func;
  assign alu_io_alu_op_alt = ID_EX_io_out_EX_alu_op_alt;
  assign alu_io_op_op1 = _T_71;
  assign alu_io_op_op2 = _T_80;
  assign dataMem_clock = clock;
  assign dataMem_io_mem_write = EX_MEM_io_out_MEM_write;
  assign dataMem_io_mem_read = EX_MEM_io_out_MEM_read;
  assign dataMem_io_mem_func = EX_MEM_io_out_MEM_func;
  assign dataMem_io_op_op1 = EX_MEM_io_out_op_op1;
  assign dataMem_io_op_op2 = EX_MEM_io_out_op_op2;
  assign fwdUnit_io_reg_w_mem = EX_MEM_io_out_WB_reg_w;
  assign fwdUnit_io_reg_w_wb = MEM_WB_io_out_WB_reg_w;
  assign fwdUnit_io_rs_rs1 = ID_EX_io_out_rs_rs1;
  assign fwdUnit_io_rs_rs2 = ID_EX_io_out_rs_rs2;
  assign fwdUnit_io_rd_mem = EX_MEM_io_out_rd;
  assign fwdUnit_io_rd_wb = MEM_WB_io_out_rd;
  assign uart_clock = clock;
  assign uart_reset = reset;
  assign uart_io_in = _GEN_1[7:0];
  assign IF_ID_clock = clock;
  assign IF_ID_io_in_pc_next = counter_io_pc_next;
  assign IF_ID_io_in_inst = instMem_io_inst;
  assign ID_EX_clock = clock;
  assign ID_EX_io_in_WB_reg_w = control_io_WB_reg_w;
  assign ID_EX_io_in_WB_rd_mem = control_io_WB_rd_mem;
  assign ID_EX_io_in_MEM_write = control_io_MEM_write;
  assign ID_EX_io_in_MEM_read = control_io_MEM_read;
  assign ID_EX_io_in_MEM_func = control_io_MEM_func;
  assign ID_EX_io_in_EX_opcode = control_io_EX_opcode;
  assign ID_EX_io_in_EX_alu_sel = control_io_EX_alu_sel;
  assign ID_EX_io_in_EX_dst_sel = control_io_EX_dst_sel;
  assign ID_EX_io_in_EX_alu_op_func = control_io_EX_alu_op_func;
  assign ID_EX_io_in_EX_alu_op_alt = control_io_EX_alu_op_alt;
  assign ID_EX_io_in_op_op1 = regs_io_op_op1;
  assign ID_EX_io_in_op_op2 = regs_io_op_op2;
  assign ID_EX_io_in_rs_rs1 = decoder_io_rs_rs1;
  assign ID_EX_io_in_rs_rs2 = decoder_io_rs_rs2;
  assign ID_EX_io_in_rd = decoder_io_rd;
  assign ID_EX_io_in_imm = decoder_io_imm;
  assign ID_EX_io_in_pc_next = IF_ID_io_out_pc_next;
  assign EX_MEM_clock = clock;
  assign EX_MEM_io_in_WB_reg_w = ID_EX_io_out_WB_reg_w;
  assign EX_MEM_io_in_WB_rd_mem = ID_EX_io_out_WB_rd_mem;
  assign EX_MEM_io_in_MEM_write = ID_EX_io_out_MEM_write;
  assign EX_MEM_io_in_MEM_read = ID_EX_io_out_MEM_read;
  assign EX_MEM_io_in_MEM_func = ID_EX_io_out_MEM_func;
  assign EX_MEM_io_in_op_op1 = alu_io_res;
  assign EX_MEM_io_in_op_op2 = ID_EX_io_out_op_op2;
  assign EX_MEM_io_in_rd = _T_81;
  assign EX_MEM_io_in_pc_next = ID_EX_io_out_pc_next;
  assign MEM_WB_clock = clock;
  assign MEM_WB_io_in_WB_reg_w = EX_MEM_io_out_WB_reg_w;
  assign MEM_WB_io_in_WB_rd_mem = EX_MEM_io_out_WB_rd_mem;
  assign MEM_WB_io_in_alu_res = EX_MEM_io_out_op_op1;
  assign MEM_WB_io_in_mem_res = dataMem_io_res;
  assign MEM_WB_io_in_rd = EX_MEM_io_out_rd;
  assign _T_51 = regs_io_op_op1 == regs_io_op_op2;
  assign _T_52 = control_io_MEM_branch & _T_51;
  assign _T_54 = uart_io_valid == 1'h0;
  assign _T_55 = _T_52 | _T_54;
  assign _T_56 = IF_ID_io_out_pc_next + decoder_io_imm;
  assign _T_57 = _T_56[31:0];
  assign _T_59 = EX_MEM_io_out_pc_next - 32'h1;
  assign _T_60 = $unsigned(_T_59);
  assign _T_61 = _T_60[31:0];
  assign _T_62 = uart_io_valid ? _T_57 : _T_61;
  assign _T_63 = uart_io_valid ? decoder_io_ctrl_opcode : 7'h0;
  assign _T_64 = uart_io_valid ? decoder_io_ctrl_funct3 : 3'h0;
  assign _T_65 = uart_io_valid ? decoder_io_ctrl_funct7 : 7'h0;
  assign _T_66 = 2'h0 == fwdUnit_io_fwd_rs1;
  assign _T_67 = _T_66 ? ID_EX_io_out_op_op1 : 32'h0;
  assign _T_68 = 2'h1 == fwdUnit_io_fwd_rs1;
  assign _T_69 = _T_68 ? regs_io_res : _T_67;
  assign _T_70 = 2'h2 == fwdUnit_io_fwd_rs1;
  assign _T_71 = _T_70 ? EX_MEM_io_out_op_op1 : _T_69;
  assign _T_72 = ID_EX_io_out_EX_alu_sel ? ID_EX_io_out_imm : EX_MEM_io_out_op_op1;
  assign _T_73 = ID_EX_io_out_EX_alu_sel ? ID_EX_io_out_imm : regs_io_res;
  assign _T_74 = ID_EX_io_out_EX_alu_sel ? ID_EX_io_out_imm : ID_EX_io_out_op_op2;
  assign _T_75 = 2'h0 == fwdUnit_io_fwd_rs2;
  assign _T_76 = _T_75 ? _T_74 : 32'h0;
  assign _T_77 = 2'h1 == fwdUnit_io_fwd_rs2;
  assign _T_78 = _T_77 ? _T_73 : _T_76;
  assign _T_79 = 2'h2 == fwdUnit_io_fwd_rs2;
  assign _T_80 = _T_79 ? _T_72 : _T_78;
  assign _T_81 = ID_EX_io_out_EX_dst_sel ? ID_EX_io_out_rd : ID_EX_io_out_rs_rs2;
  assign _T_82 = MEM_WB_io_out_WB_rd_mem ? MEM_WB_io_out_mem_res : MEM_WB_io_out_alu_res;
  assign _T_84 = dataMem_io_op_op1 == 32'h401;
  assign _T_85 = EX_MEM_io_out_MEM_write & _T_84;
  assign _GEN_0 = dataMem_io_op_op2;
  assign _T_87 = _T_85 == 1'h0;
  assign _GEN_1 = _T_87 ? 32'h0 : _GEN_0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_6 = {1{$random}};
  _GEN_2 = _GEN_6[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_7 = {1{$random}};
  _GEN_3 = _GEN_7[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_8 = {1{$random}};
  _GEN_4 = _GEN_8[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  _GEN_9 = {1{$random}};
  _GEN_5 = _GEN_9[0:0];
  `endif
  end
`endif
endmodule
